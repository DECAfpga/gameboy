
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"54",x"7c",x"38",x"00"),
     1 => (x"00",x"18",x"5c",x"54"),
     2 => (x"7f",x"7e",x"04",x"00"),
     3 => (x"00",x"00",x"05",x"05"),
     4 => (x"a4",x"bc",x"18",x"00"),
     5 => (x"00",x"7c",x"fc",x"a4"),
     6 => (x"04",x"7f",x"7f",x"00"),
     7 => (x"00",x"78",x"7c",x"04"),
     8 => (x"3d",x"00",x"00",x"00"),
     9 => (x"00",x"00",x"40",x"7d"),
    10 => (x"80",x"80",x"80",x"00"),
    11 => (x"00",x"00",x"7d",x"fd"),
    12 => (x"10",x"7f",x"7f",x"00"),
    13 => (x"00",x"44",x"6c",x"38"),
    14 => (x"3f",x"00",x"00",x"00"),
    15 => (x"00",x"00",x"40",x"7f"),
    16 => (x"18",x"0c",x"7c",x"7c"),
    17 => (x"00",x"78",x"7c",x"0c"),
    18 => (x"04",x"7c",x"7c",x"00"),
    19 => (x"00",x"78",x"7c",x"04"),
    20 => (x"44",x"7c",x"38",x"00"),
    21 => (x"00",x"38",x"7c",x"44"),
    22 => (x"24",x"fc",x"fc",x"00"),
    23 => (x"00",x"18",x"3c",x"24"),
    24 => (x"24",x"3c",x"18",x"00"),
    25 => (x"00",x"fc",x"fc",x"24"),
    26 => (x"04",x"7c",x"7c",x"00"),
    27 => (x"00",x"08",x"0c",x"04"),
    28 => (x"54",x"5c",x"48",x"00"),
    29 => (x"00",x"20",x"74",x"54"),
    30 => (x"7f",x"3f",x"04",x"00"),
    31 => (x"00",x"00",x"44",x"44"),
    32 => (x"40",x"7c",x"3c",x"00"),
    33 => (x"00",x"7c",x"7c",x"40"),
    34 => (x"60",x"3c",x"1c",x"00"),
    35 => (x"00",x"1c",x"3c",x"60"),
    36 => (x"30",x"60",x"7c",x"3c"),
    37 => (x"00",x"3c",x"7c",x"60"),
    38 => (x"10",x"38",x"6c",x"44"),
    39 => (x"00",x"44",x"6c",x"38"),
    40 => (x"e0",x"bc",x"1c",x"00"),
    41 => (x"00",x"1c",x"3c",x"60"),
    42 => (x"74",x"64",x"44",x"00"),
    43 => (x"00",x"44",x"4c",x"5c"),
    44 => (x"3e",x"08",x"08",x"00"),
    45 => (x"00",x"41",x"41",x"77"),
    46 => (x"7f",x"00",x"00",x"00"),
    47 => (x"00",x"00",x"00",x"7f"),
    48 => (x"77",x"41",x"41",x"00"),
    49 => (x"00",x"08",x"08",x"3e"),
    50 => (x"03",x"01",x"01",x"02"),
    51 => (x"00",x"01",x"02",x"02"),
    52 => (x"7f",x"7f",x"7f",x"7f"),
    53 => (x"00",x"7f",x"7f",x"7f"),
    54 => (x"1c",x"1c",x"08",x"08"),
    55 => (x"7f",x"7f",x"3e",x"3e"),
    56 => (x"3e",x"3e",x"7f",x"7f"),
    57 => (x"08",x"08",x"1c",x"1c"),
    58 => (x"7c",x"18",x"10",x"00"),
    59 => (x"00",x"10",x"18",x"7c"),
    60 => (x"7c",x"30",x"10",x"00"),
    61 => (x"00",x"10",x"30",x"7c"),
    62 => (x"60",x"60",x"30",x"10"),
    63 => (x"00",x"06",x"1e",x"78"),
    64 => (x"18",x"3c",x"66",x"42"),
    65 => (x"00",x"42",x"66",x"3c"),
    66 => (x"c2",x"6a",x"38",x"78"),
    67 => (x"00",x"38",x"6c",x"c6"),
    68 => (x"60",x"00",x"00",x"60"),
    69 => (x"00",x"60",x"00",x"00"),
    70 => (x"5c",x"5b",x"5e",x"0e"),
    71 => (x"86",x"fc",x"0e",x"5d"),
    72 => (x"e8",x"c2",x"7e",x"71"),
    73 => (x"c0",x"4c",x"bf",x"e8"),
    74 => (x"c4",x"1e",x"c0",x"4b"),
    75 => (x"c4",x"02",x"ab",x"66"),
    76 => (x"c2",x"4d",x"c0",x"87"),
    77 => (x"75",x"4d",x"c1",x"87"),
    78 => (x"ee",x"49",x"73",x"1e"),
    79 => (x"86",x"c8",x"87",x"e2"),
    80 => (x"ef",x"49",x"e0",x"c0"),
    81 => (x"a4",x"c4",x"87",x"eb"),
    82 => (x"f0",x"49",x"6a",x"4a"),
    83 => (x"c9",x"f1",x"87",x"f2"),
    84 => (x"c1",x"84",x"cc",x"87"),
    85 => (x"ab",x"b7",x"c8",x"83"),
    86 => (x"87",x"cd",x"ff",x"04"),
    87 => (x"4d",x"26",x"8e",x"fc"),
    88 => (x"4b",x"26",x"4c",x"26"),
    89 => (x"71",x"1e",x"4f",x"26"),
    90 => (x"ec",x"e8",x"c2",x"4a"),
    91 => (x"ec",x"e8",x"c2",x"5a"),
    92 => (x"49",x"78",x"c7",x"48"),
    93 => (x"26",x"87",x"e1",x"fe"),
    94 => (x"1e",x"73",x"1e",x"4f"),
    95 => (x"b7",x"c0",x"4a",x"71"),
    96 => (x"87",x"d3",x"03",x"aa"),
    97 => (x"bf",x"f4",x"d4",x"c2"),
    98 => (x"c1",x"87",x"c4",x"05"),
    99 => (x"c0",x"87",x"c2",x"4b"),
   100 => (x"f8",x"d4",x"c2",x"4b"),
   101 => (x"c2",x"87",x"c4",x"5b"),
   102 => (x"fc",x"5a",x"f8",x"d4"),
   103 => (x"f4",x"d4",x"c2",x"48"),
   104 => (x"c1",x"4a",x"78",x"bf"),
   105 => (x"a2",x"c0",x"c1",x"9a"),
   106 => (x"87",x"e7",x"ec",x"49"),
   107 => (x"4f",x"26",x"4b",x"26"),
   108 => (x"c4",x"4a",x"71",x"1e"),
   109 => (x"49",x"72",x"1e",x"66"),
   110 => (x"fc",x"87",x"f1",x"eb"),
   111 => (x"1e",x"4f",x"26",x"8e"),
   112 => (x"c3",x"48",x"d4",x"ff"),
   113 => (x"d0",x"ff",x"78",x"ff"),
   114 => (x"78",x"e1",x"c0",x"48"),
   115 => (x"c1",x"48",x"d4",x"ff"),
   116 => (x"c4",x"48",x"71",x"78"),
   117 => (x"08",x"d4",x"ff",x"30"),
   118 => (x"48",x"d0",x"ff",x"78"),
   119 => (x"26",x"78",x"e0",x"c0"),
   120 => (x"5b",x"5e",x"0e",x"4f"),
   121 => (x"f0",x"0e",x"5d",x"5c"),
   122 => (x"48",x"a6",x"c8",x"86"),
   123 => (x"bf",x"ec",x"78",x"c0"),
   124 => (x"c2",x"80",x"fc",x"7e"),
   125 => (x"78",x"bf",x"e8",x"e8"),
   126 => (x"bf",x"f0",x"e8",x"c2"),
   127 => (x"4c",x"bf",x"e8",x"4d"),
   128 => (x"bf",x"f4",x"d4",x"c2"),
   129 => (x"87",x"f9",x"e3",x"49"),
   130 => (x"f6",x"e8",x"49",x"c7"),
   131 => (x"c2",x"49",x"70",x"87"),
   132 => (x"87",x"cf",x"05",x"99"),
   133 => (x"bf",x"ec",x"d4",x"c2"),
   134 => (x"6e",x"b9",x"ff",x"49"),
   135 => (x"02",x"99",x"c1",x"99"),
   136 => (x"cb",x"87",x"c0",x"c2"),
   137 => (x"cf",x"cc",x"49",x"ee"),
   138 => (x"58",x"a6",x"d0",x"87"),
   139 => (x"d2",x"e8",x"49",x"c7"),
   140 => (x"05",x"98",x"70",x"87"),
   141 => (x"49",x"6e",x"87",x"c8"),
   142 => (x"c1",x"02",x"99",x"c1"),
   143 => (x"66",x"cc",x"87",x"c2"),
   144 => (x"7e",x"bf",x"ec",x"4b"),
   145 => (x"bf",x"f4",x"d4",x"c2"),
   146 => (x"87",x"f5",x"e2",x"49"),
   147 => (x"f3",x"cb",x"49",x"73"),
   148 => (x"02",x"98",x"70",x"87"),
   149 => (x"d4",x"c2",x"87",x"d7"),
   150 => (x"c1",x"49",x"bf",x"d4"),
   151 => (x"d8",x"d4",x"c2",x"b9"),
   152 => (x"da",x"fd",x"71",x"59"),
   153 => (x"49",x"ee",x"cb",x"87"),
   154 => (x"70",x"87",x"cd",x"cb"),
   155 => (x"e7",x"49",x"c7",x"4b"),
   156 => (x"98",x"70",x"87",x"d1"),
   157 => (x"87",x"c9",x"ff",x"05"),
   158 => (x"99",x"c1",x"49",x"6e"),
   159 => (x"87",x"c1",x"ff",x"05"),
   160 => (x"bf",x"f4",x"d4",x"c2"),
   161 => (x"c2",x"ba",x"c1",x"4a"),
   162 => (x"fc",x"5a",x"f8",x"d4"),
   163 => (x"c1",x"0a",x"7a",x"0a"),
   164 => (x"a2",x"c0",x"c1",x"9a"),
   165 => (x"87",x"fb",x"e8",x"49"),
   166 => (x"e6",x"49",x"da",x"c1"),
   167 => (x"a6",x"c8",x"87",x"e5"),
   168 => (x"c2",x"78",x"c1",x"48"),
   169 => (x"6e",x"48",x"ec",x"d4"),
   170 => (x"f4",x"d4",x"c2",x"78"),
   171 => (x"c7",x"c1",x"05",x"bf"),
   172 => (x"c0",x"c0",x"c8",x"87"),
   173 => (x"e0",x"d5",x"c2",x"4b"),
   174 => (x"49",x"15",x"4d",x"7e"),
   175 => (x"87",x"c3",x"e6",x"49"),
   176 => (x"c0",x"02",x"98",x"70"),
   177 => (x"b4",x"73",x"87",x"c2"),
   178 => (x"05",x"2b",x"b7",x"c1"),
   179 => (x"74",x"87",x"eb",x"ff"),
   180 => (x"99",x"ff",x"c3",x"49"),
   181 => (x"49",x"c0",x"1e",x"71"),
   182 => (x"74",x"87",x"d5",x"fb"),
   183 => (x"29",x"b7",x"c8",x"49"),
   184 => (x"49",x"c1",x"1e",x"71"),
   185 => (x"c8",x"87",x"c9",x"fb"),
   186 => (x"49",x"fd",x"c3",x"86"),
   187 => (x"c3",x"87",x"d4",x"e5"),
   188 => (x"ce",x"e5",x"49",x"fa"),
   189 => (x"87",x"d1",x"c8",x"87"),
   190 => (x"ff",x"c3",x"49",x"74"),
   191 => (x"2c",x"b7",x"c8",x"99"),
   192 => (x"9c",x"74",x"b4",x"71"),
   193 => (x"ff",x"87",x"df",x"02"),
   194 => (x"49",x"7e",x"bf",x"c8"),
   195 => (x"bf",x"f0",x"d4",x"c2"),
   196 => (x"a9",x"e0",x"c2",x"89"),
   197 => (x"87",x"c5",x"c0",x"03"),
   198 => (x"cf",x"c0",x"4c",x"c0"),
   199 => (x"f0",x"d4",x"c2",x"87"),
   200 => (x"c0",x"78",x"6e",x"48"),
   201 => (x"d4",x"c2",x"87",x"c6"),
   202 => (x"78",x"c0",x"48",x"f0"),
   203 => (x"99",x"c8",x"49",x"74"),
   204 => (x"87",x"ce",x"c0",x"05"),
   205 => (x"e4",x"49",x"f5",x"c3"),
   206 => (x"49",x"70",x"87",x"c9"),
   207 => (x"c0",x"02",x"99",x"c2"),
   208 => (x"e8",x"c2",x"87",x"ea"),
   209 => (x"c0",x"02",x"bf",x"ec"),
   210 => (x"c1",x"48",x"87",x"ca"),
   211 => (x"f0",x"e8",x"c2",x"88"),
   212 => (x"87",x"d3",x"c0",x"58"),
   213 => (x"c1",x"48",x"66",x"c4"),
   214 => (x"7e",x"70",x"80",x"e0"),
   215 => (x"c0",x"02",x"bf",x"6e"),
   216 => (x"ff",x"4b",x"87",x"c5"),
   217 => (x"c8",x"0f",x"73",x"49"),
   218 => (x"78",x"c1",x"48",x"a6"),
   219 => (x"99",x"c4",x"49",x"74"),
   220 => (x"87",x"ce",x"c0",x"05"),
   221 => (x"e3",x"49",x"f2",x"c3"),
   222 => (x"49",x"70",x"87",x"c9"),
   223 => (x"c0",x"02",x"99",x"c2"),
   224 => (x"e8",x"c2",x"87",x"f0"),
   225 => (x"48",x"7e",x"bf",x"ec"),
   226 => (x"03",x"a8",x"b7",x"c7"),
   227 => (x"6e",x"87",x"cb",x"c0"),
   228 => (x"c2",x"80",x"c1",x"48"),
   229 => (x"c0",x"58",x"f0",x"e8"),
   230 => (x"66",x"c4",x"87",x"d3"),
   231 => (x"80",x"e0",x"c1",x"48"),
   232 => (x"bf",x"6e",x"7e",x"70"),
   233 => (x"87",x"c5",x"c0",x"02"),
   234 => (x"73",x"49",x"fe",x"4b"),
   235 => (x"48",x"a6",x"c8",x"0f"),
   236 => (x"fd",x"c3",x"78",x"c1"),
   237 => (x"87",x"cb",x"e2",x"49"),
   238 => (x"99",x"c2",x"49",x"70"),
   239 => (x"87",x"e6",x"c0",x"02"),
   240 => (x"bf",x"ec",x"e8",x"c2"),
   241 => (x"87",x"c9",x"c0",x"02"),
   242 => (x"48",x"ec",x"e8",x"c2"),
   243 => (x"d0",x"c0",x"78",x"c0"),
   244 => (x"4a",x"66",x"c4",x"87"),
   245 => (x"6a",x"82",x"e0",x"c1"),
   246 => (x"87",x"c5",x"c0",x"02"),
   247 => (x"73",x"49",x"fd",x"4b"),
   248 => (x"48",x"a6",x"c8",x"0f"),
   249 => (x"fa",x"c3",x"78",x"c1"),
   250 => (x"87",x"d7",x"e1",x"49"),
   251 => (x"99",x"c2",x"49",x"70"),
   252 => (x"87",x"ed",x"c0",x"02"),
   253 => (x"bf",x"ec",x"e8",x"c2"),
   254 => (x"a8",x"b7",x"c7",x"48"),
   255 => (x"87",x"c9",x"c0",x"03"),
   256 => (x"48",x"ec",x"e8",x"c2"),
   257 => (x"d3",x"c0",x"78",x"c7"),
   258 => (x"48",x"66",x"c4",x"87"),
   259 => (x"70",x"80",x"e0",x"c1"),
   260 => (x"02",x"bf",x"6e",x"7e"),
   261 => (x"4b",x"87",x"c5",x"c0"),
   262 => (x"0f",x"73",x"49",x"fc"),
   263 => (x"c1",x"48",x"a6",x"c8"),
   264 => (x"c3",x"48",x"74",x"78"),
   265 => (x"7e",x"70",x"98",x"f0"),
   266 => (x"c0",x"05",x"98",x"48"),
   267 => (x"da",x"c1",x"87",x"ce"),
   268 => (x"87",x"cf",x"e0",x"49"),
   269 => (x"99",x"c2",x"49",x"70"),
   270 => (x"87",x"d0",x"c2",x"02"),
   271 => (x"c3",x"49",x"ee",x"cb"),
   272 => (x"a6",x"d0",x"87",x"f6"),
   273 => (x"e4",x"e8",x"c2",x"58"),
   274 => (x"c2",x"50",x"c0",x"48"),
   275 => (x"bf",x"97",x"e4",x"e8"),
   276 => (x"87",x"d8",x"c1",x"05"),
   277 => (x"cd",x"c0",x"05",x"6e"),
   278 => (x"49",x"da",x"c1",x"87"),
   279 => (x"87",x"e3",x"df",x"ff"),
   280 => (x"c1",x"02",x"98",x"70"),
   281 => (x"bf",x"e8",x"87",x"c6"),
   282 => (x"ff",x"c3",x"49",x"4b"),
   283 => (x"2b",x"b7",x"c8",x"99"),
   284 => (x"d4",x"c2",x"b3",x"71"),
   285 => (x"ff",x"49",x"bf",x"f4"),
   286 => (x"cc",x"87",x"c6",x"da"),
   287 => (x"c3",x"c3",x"49",x"66"),
   288 => (x"02",x"98",x"70",x"87"),
   289 => (x"c2",x"87",x"c6",x"c0"),
   290 => (x"c1",x"48",x"e4",x"e8"),
   291 => (x"e4",x"e8",x"c2",x"50"),
   292 => (x"c0",x"05",x"bf",x"97"),
   293 => (x"49",x"73",x"87",x"d6"),
   294 => (x"05",x"99",x"f0",x"c3"),
   295 => (x"c1",x"87",x"c7",x"ff"),
   296 => (x"de",x"ff",x"49",x"da"),
   297 => (x"98",x"70",x"87",x"dd"),
   298 => (x"87",x"fa",x"fe",x"05"),
   299 => (x"c2",x"48",x"a6",x"cc"),
   300 => (x"78",x"bf",x"ec",x"e8"),
   301 => (x"cc",x"49",x"66",x"cc"),
   302 => (x"48",x"66",x"c4",x"91"),
   303 => (x"7e",x"70",x"80",x"71"),
   304 => (x"c0",x"02",x"bf",x"6e"),
   305 => (x"cc",x"4b",x"87",x"c6"),
   306 => (x"0f",x"73",x"49",x"66"),
   307 => (x"c0",x"02",x"9d",x"75"),
   308 => (x"02",x"6d",x"87",x"e9"),
   309 => (x"6d",x"87",x"e4",x"c0"),
   310 => (x"e6",x"dd",x"ff",x"49"),
   311 => (x"c1",x"49",x"70",x"87"),
   312 => (x"cb",x"c0",x"02",x"99"),
   313 => (x"4b",x"a5",x"c4",x"87"),
   314 => (x"bf",x"ec",x"e8",x"c2"),
   315 => (x"0f",x"4b",x"6b",x"49"),
   316 => (x"c0",x"02",x"85",x"c8"),
   317 => (x"05",x"6d",x"87",x"c5"),
   318 => (x"c8",x"87",x"dc",x"ff"),
   319 => (x"c8",x"c0",x"02",x"66"),
   320 => (x"ec",x"e8",x"c2",x"87"),
   321 => (x"cf",x"f0",x"49",x"bf"),
   322 => (x"26",x"8e",x"f0",x"87"),
   323 => (x"26",x"4c",x"26",x"4d"),
   324 => (x"00",x"4f",x"26",x"4b"),
   325 => (x"00",x"00",x"00",x"00"),
   326 => (x"00",x"00",x"00",x"10"),
   327 => (x"14",x"11",x"12",x"58"),
   328 => (x"23",x"1c",x"1b",x"1d"),
   329 => (x"94",x"91",x"59",x"5a"),
   330 => (x"f4",x"eb",x"f2",x"f5"),
   331 => (x"00",x"00",x"00",x"00"),
   332 => (x"00",x"00",x"00",x"00"),
   333 => (x"00",x"00",x"00",x"00"),
   334 => (x"ff",x"4a",x"71",x"1e"),
   335 => (x"72",x"49",x"bf",x"c8"),
   336 => (x"4f",x"26",x"48",x"a1"),
   337 => (x"bf",x"c8",x"ff",x"1e"),
   338 => (x"c0",x"c0",x"fe",x"89"),
   339 => (x"a9",x"c0",x"c0",x"c0"),
   340 => (x"c0",x"87",x"c4",x"01"),
   341 => (x"c1",x"87",x"c2",x"4a"),
   342 => (x"26",x"48",x"72",x"4a"),
   343 => (x"00",x"00",x"00",x"4f"),
   344 => (x"11",x"14",x"12",x"58"),
   345 => (x"23",x"1c",x"1b",x"1d"),
   346 => (x"91",x"94",x"59",x"5a"),
   347 => (x"f4",x"eb",x"f2",x"f5"),
   348 => (x"00",x"00",x"25",x"74"),
   349 => (x"4f",x"54",x"55",x"41"),
   350 => (x"54",x"4f",x"4f",x"42"),
   351 => (x"17",x"00",x"42",x"47"),
   352 => (x"17",x"00",x"00",x"1a"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

