library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"d4eac287",
    12 => x"48c0c84e",
    13 => x"d5c128c2",
    14 => x"ead6e5ea",
    15 => x"c1467149",
    16 => x"87f90188",
    17 => x"49d4eac2",
    18 => x"48e4d7c2",
    19 => x"0389d089",
    20 => x"404040c0",
    21 => x"d087f640",
    22 => x"50c00581",
    23 => x"f90589c1",
    24 => x"e4d7c287",
    25 => x"e0d7c24d",
    26 => x"02ad744c",
    27 => x"0f2487c4",
    28 => x"e2c187f7",
    29 => x"d7c287d4",
    30 => x"d7c24de4",
    31 => x"ad744ce4",
    32 => x"c487c602",
    33 => x"f50f6c8c",
    34 => x"87fd0087",
    35 => x"7186fc1e",
    36 => x"49c0ff4a",
    37 => x"c0c44869",
    38 => x"487e7098",
    39 => x"87f40298",
    40 => x"fc487972",
    41 => x"0e4f268e",
    42 => x"0e5c5b5e",
    43 => x"4cc04b71",
    44 => x"029a4a13",
    45 => x"497287cd",
    46 => x"c187d1ff",
    47 => x"9a4a1384",
    48 => x"7487f305",
    49 => x"264c2648",
    50 => x"1e4f264b",
    51 => x"1e731e72",
    52 => x"02114812",
    53 => x"c34b87ca",
    54 => x"739b98df",
    55 => x"87f00288",
    56 => x"4a264b26",
    57 => x"731e4f26",
    58 => x"c11e721e",
    59 => x"87ca048b",
    60 => x"02114812",
    61 => x"028887c4",
    62 => x"4a2687f1",
    63 => x"4f264b26",
    64 => x"731e741e",
    65 => x"c11e721e",
    66 => x"87cf048b",
    67 => x"02114812",
    68 => x"df4c87c9",
    69 => x"88749c98",
    70 => x"2687ec02",
    71 => x"264b264a",
    72 => x"1e4f264c",
    73 => x"73814873",
    74 => x"87c502a9",
    75 => x"f6055312",
    76 => x"0e4f2687",
    77 => x"0e5c5b5e",
    78 => x"d4ff4a71",
    79 => x"4b66cc4c",
    80 => x"718bc149",
    81 => x"87ce0299",
    82 => x"6c7cffc3",
    83 => x"c1497352",
    84 => x"0599718b",
    85 => x"4c2687f2",
    86 => x"4f264b26",
    87 => x"ff1e731e",
    88 => x"ffc34bd4",
    89 => x"c34a6b7b",
    90 => x"496b7bff",
    91 => x"b17232c8",
    92 => x"6b7bffc3",
    93 => x"7131c84a",
    94 => x"7bffc3b2",
    95 => x"32c8496b",
    96 => x"4871b172",
    97 => x"4f264b26",
    98 => x"5c5b5e0e",
    99 => x"4d710e5d",
   100 => x"754cd4ff",
   101 => x"98ffc348",
   102 => x"d7c27c70",
   103 => x"c805bfe4",
   104 => x"4866d087",
   105 => x"a6d430c9",
   106 => x"4966d058",
   107 => x"487129d8",
   108 => x"7098ffc3",
   109 => x"4966d07c",
   110 => x"487129d0",
   111 => x"7098ffc3",
   112 => x"4966d07c",
   113 => x"487129c8",
   114 => x"7098ffc3",
   115 => x"4866d07c",
   116 => x"7098ffc3",
   117 => x"d049757c",
   118 => x"c3487129",
   119 => x"7c7098ff",
   120 => x"f0c94b6c",
   121 => x"ffc34aff",
   122 => x"87cf05ab",
   123 => x"6c7c7149",
   124 => x"028ac14b",
   125 => x"ab7187c5",
   126 => x"7387f202",
   127 => x"264d2648",
   128 => x"264b264c",
   129 => x"49c01e4f",
   130 => x"c348d4ff",
   131 => x"81c178ff",
   132 => x"a9b7c8c3",
   133 => x"2687f104",
   134 => x"5b5e0e4f",
   135 => x"c00e5d5c",
   136 => x"f7c1f0ff",
   137 => x"c0c0c14d",
   138 => x"4bc0c0c0",
   139 => x"c487d6ff",
   140 => x"c04cdff8",
   141 => x"fd49751e",
   142 => x"86c487ce",
   143 => x"c005a8c1",
   144 => x"d4ff87e5",
   145 => x"78ffc348",
   146 => x"e1c01e73",
   147 => x"49e9c1f0",
   148 => x"c487f5fc",
   149 => x"05987086",
   150 => x"d4ff87ca",
   151 => x"78ffc348",
   152 => x"87cb48c1",
   153 => x"c187defe",
   154 => x"c6ff058c",
   155 => x"2648c087",
   156 => x"264c264d",
   157 => x"0e4f264b",
   158 => x"0e5c5b5e",
   159 => x"c1f0ffc0",
   160 => x"d4ff4cc1",
   161 => x"78ffc348",
   162 => x"f849fcca",
   163 => x"4bd387d9",
   164 => x"49741ec0",
   165 => x"c487f1fb",
   166 => x"05987086",
   167 => x"d4ff87ca",
   168 => x"78ffc348",
   169 => x"87cb48c1",
   170 => x"c187dafd",
   171 => x"dfff058b",
   172 => x"2648c087",
   173 => x"264b264c",
   174 => x"0000004f",
   175 => x"00444d43",
   176 => x"43484453",
   177 => x"69616620",
   178 => x"000a216c",
   179 => x"52524549",
   180 => x"00000000",
   181 => x"00495053",
   182 => x"74697257",
   183 => x"61662065",
   184 => x"64656c69",
   185 => x"5e0e000a",
   186 => x"0e5d5c5b",
   187 => x"ff4dffc3",
   188 => x"d0fc4bd4",
   189 => x"1eeac687",
   190 => x"c1f0e1c0",
   191 => x"c7fa49c8",
   192 => x"c186c487",
   193 => x"87c802a8",
   194 => x"c087ecfd",
   195 => x"87e8c148",
   196 => x"7087c9f9",
   197 => x"ffffcf49",
   198 => x"a9eac699",
   199 => x"fd87c802",
   200 => x"48c087d5",
   201 => x"7587d1c1",
   202 => x"4cf1c07b",
   203 => x"7087eafb",
   204 => x"ecc00298",
   205 => x"c01ec087",
   206 => x"fac1f0ff",
   207 => x"87c8f949",
   208 => x"987086c4",
   209 => x"7587da05",
   210 => x"75496b7b",
   211 => x"757b757b",
   212 => x"c17b757b",
   213 => x"c40299c0",
   214 => x"db48c187",
   215 => x"d748c087",
   216 => x"05acc287",
   217 => x"c0cb87ca",
   218 => x"87fbf449",
   219 => x"87c848c0",
   220 => x"fe058cc1",
   221 => x"48c087f6",
   222 => x"4c264d26",
   223 => x"4f264b26",
   224 => x"5c5b5e0e",
   225 => x"d0ff0e5d",
   226 => x"d0e5c04d",
   227 => x"c24cc0c1",
   228 => x"c148e4d7",
   229 => x"49d4cb78",
   230 => x"c787ccf4",
   231 => x"f97dc24b",
   232 => x"7dc387e3",
   233 => x"49741ec0",
   234 => x"c487ddf7",
   235 => x"05a8c186",
   236 => x"c24b87c1",
   237 => x"87cb05ab",
   238 => x"f349cccb",
   239 => x"48c087e9",
   240 => x"c187f6c0",
   241 => x"d4ff058b",
   242 => x"87dafc87",
   243 => x"58e8d7c2",
   244 => x"cd059870",
   245 => x"c01ec187",
   246 => x"d0c1f0ff",
   247 => x"87e8f649",
   248 => x"d4ff86c4",
   249 => x"78ffc348",
   250 => x"c287c3c3",
   251 => x"c258ecd7",
   252 => x"48d4ff7d",
   253 => x"c178ffc3",
   254 => x"264d2648",
   255 => x"264b264c",
   256 => x"5b5e0e4f",
   257 => x"fc0e5d5c",
   258 => x"ff4b7186",
   259 => x"7ec04cd4",
   260 => x"dfcdeec5",
   261 => x"7cffc34a",
   262 => x"fec3486c",
   263 => x"f8c005a8",
   264 => x"734d7487",
   265 => x"87cc029b",
   266 => x"731e66d4",
   267 => x"87c3f449",
   268 => x"87d486c4",
   269 => x"c448d0ff",
   270 => x"66d478d1",
   271 => x"7dffc34a",
   272 => x"f8058ac1",
   273 => x"5aa6d887",
   274 => x"7c7cffc3",
   275 => x"c5059b73",
   276 => x"48d0ff87",
   277 => x"4ac178d0",
   278 => x"058ac17e",
   279 => x"6e87f6fe",
   280 => x"268efc48",
   281 => x"264c264d",
   282 => x"1e4f264b",
   283 => x"4a711e73",
   284 => x"d4ff4bc0",
   285 => x"78ffc348",
   286 => x"c448d0ff",
   287 => x"d4ff78c3",
   288 => x"78ffc348",
   289 => x"ffc01e72",
   290 => x"49d1c1f0",
   291 => x"c487f9f3",
   292 => x"05987086",
   293 => x"c0c887d2",
   294 => x"4966cc1e",
   295 => x"c487e2fd",
   296 => x"ff4b7086",
   297 => x"78c248d0",
   298 => x"4b264873",
   299 => x"5e0e4f26",
   300 => x"0e5d5c5b",
   301 => x"ffc01ec0",
   302 => x"49c9c1f0",
   303 => x"d287c9f3",
   304 => x"f4d7c21e",
   305 => x"87f9fc49",
   306 => x"4cc086c8",
   307 => x"b7d284c1",
   308 => x"87f804ac",
   309 => x"97f4d7c2",
   310 => x"c0c349bf",
   311 => x"a9c0c199",
   312 => x"87e7c005",
   313 => x"97fbd7c2",
   314 => x"31d049bf",
   315 => x"97fcd7c2",
   316 => x"32c84abf",
   317 => x"d7c2b172",
   318 => x"4abf97fd",
   319 => x"cf4c71b1",
   320 => x"9cffffff",
   321 => x"34ca84c1",
   322 => x"c287e7c1",
   323 => x"bf97fdd7",
   324 => x"c631c149",
   325 => x"fed7c299",
   326 => x"c74abf97",
   327 => x"b1722ab7",
   328 => x"97f9d7c2",
   329 => x"cf4d4abf",
   330 => x"fad7c29d",
   331 => x"c34abf97",
   332 => x"c232ca9a",
   333 => x"bf97fbd7",
   334 => x"7333c24b",
   335 => x"fcd7c2b2",
   336 => x"c34bbf97",
   337 => x"b7c69bc0",
   338 => x"c2b2732b",
   339 => x"7148c181",
   340 => x"c1497030",
   341 => x"70307548",
   342 => x"c14c724d",
   343 => x"c8947184",
   344 => x"06adb7c0",
   345 => x"34c187cc",
   346 => x"c0c82db7",
   347 => x"ff01adb7",
   348 => x"487487f4",
   349 => x"4c264d26",
   350 => x"4f264b26",
   351 => x"5c5b5e0e",
   352 => x"86f80e5d",
   353 => x"48dce0c2",
   354 => x"d8c278c0",
   355 => x"49c01ed4",
   356 => x"c487d8fb",
   357 => x"05987086",
   358 => x"48c087c5",
   359 => x"c087f1c8",
   360 => x"c27ec14d",
   361 => x"df4acad9",
   362 => x"4bc849e8",
   363 => x"7087f7ec",
   364 => x"87c20598",
   365 => x"d9c27ec0",
   366 => x"f4df4ae6",
   367 => x"ec4bc849",
   368 => x"987087e4",
   369 => x"c087c205",
   370 => x"c0026e7e",
   371 => x"dfc287fd",
   372 => x"c24dbfda",
   373 => x"bf9fd2e0",
   374 => x"d6c5487e",
   375 => x"c705a8ea",
   376 => x"dadfc287",
   377 => x"87ce4dbf",
   378 => x"e9ca486e",
   379 => x"c502a8d5",
   380 => x"c748c087",
   381 => x"d8c287da",
   382 => x"49751ed4",
   383 => x"c487ecf9",
   384 => x"05987086",
   385 => x"48c087c5",
   386 => x"c287c5c7",
   387 => x"c04ae6d9",
   388 => x"c849c0e0",
   389 => x"87ceeb4b",
   390 => x"c8059870",
   391 => x"dce0c287",
   392 => x"d778c148",
   393 => x"cad9c287",
   394 => x"cce0c04a",
   395 => x"ea4bc849",
   396 => x"987087f4",
   397 => x"c087c502",
   398 => x"87d4c648",
   399 => x"97d2e0c2",
   400 => x"d5c149bf",
   401 => x"87cd05a9",
   402 => x"97d3e0c2",
   403 => x"eac249bf",
   404 => x"c5c002a9",
   405 => x"c548c087",
   406 => x"d8c287f6",
   407 => x"7ebf97d4",
   408 => x"a8e9c348",
   409 => x"87cec002",
   410 => x"ebc3486e",
   411 => x"c5c002a8",
   412 => x"c548c087",
   413 => x"d8c287da",
   414 => x"49bf97df",
   415 => x"ccc00599",
   416 => x"e0d8c287",
   417 => x"c249bf97",
   418 => x"c5c002a9",
   419 => x"c448c087",
   420 => x"d8c287fe",
   421 => x"48bf97e1",
   422 => x"58d8e0c2",
   423 => x"c1484c70",
   424 => x"dce0c288",
   425 => x"e2d8c258",
   426 => x"7549bf97",
   427 => x"e3d8c281",
   428 => x"c84abf97",
   429 => x"7ea17232",
   430 => x"48ece4c2",
   431 => x"d8c2786e",
   432 => x"48bf97e4",
   433 => x"c258a6c8",
   434 => x"02bfdce0",
   435 => x"c287ccc2",
   436 => x"df4ae6d9",
   437 => x"4bc849dc",
   438 => x"7087cbe8",
   439 => x"c5c00298",
   440 => x"c348c087",
   441 => x"e0c287ea",
   442 => x"c24cbfd4",
   443 => x"c25cc0e5",
   444 => x"bf97f9d8",
   445 => x"c231c849",
   446 => x"bf97f8d8",
   447 => x"c249a14a",
   448 => x"bf97fad8",
   449 => x"7232d04a",
   450 => x"d8c249a1",
   451 => x"4abf97fb",
   452 => x"a17232d8",
   453 => x"9166c449",
   454 => x"bfece4c2",
   455 => x"f4e4c281",
   456 => x"c1d9c259",
   457 => x"c84abf97",
   458 => x"c0d9c232",
   459 => x"a24bbf97",
   460 => x"c2d9c24a",
   461 => x"d04bbf97",
   462 => x"4aa27333",
   463 => x"97c3d9c2",
   464 => x"9bcf4bbf",
   465 => x"a27333d8",
   466 => x"f8e4c24a",
   467 => x"748ac25a",
   468 => x"f8e4c292",
   469 => x"78a17248",
   470 => x"c287c1c1",
   471 => x"bf97e6d8",
   472 => x"c231c849",
   473 => x"bf97e5d8",
   474 => x"c549a14a",
   475 => x"81ffc731",
   476 => x"e5c229c9",
   477 => x"d8c259c0",
   478 => x"4abf97eb",
   479 => x"d8c232c8",
   480 => x"4bbf97ea",
   481 => x"66c44aa2",
   482 => x"c2826e92",
   483 => x"c25afce4",
   484 => x"c048f4e4",
   485 => x"f0e4c278",
   486 => x"78a17248",
   487 => x"48c0e5c2",
   488 => x"bff4e4c2",
   489 => x"c4e5c278",
   490 => x"f8e4c248",
   491 => x"e0c278bf",
   492 => x"c002bfdc",
   493 => x"487487c9",
   494 => x"7e7030c4",
   495 => x"c287c9c0",
   496 => x"48bffce4",
   497 => x"7e7030c4",
   498 => x"48e0e0c2",
   499 => x"48c1786e",
   500 => x"4d268ef8",
   501 => x"4b264c26",
   502 => x"00004f26",
   503 => x"33544146",
   504 => x"20202032",
   505 => x"00000000",
   506 => x"31544146",
   507 => x"20202036",
   508 => x"00000000",
   509 => x"33544146",
   510 => x"20202032",
   511 => x"00000000",
   512 => x"33544146",
   513 => x"20202032",
   514 => x"00000000",
   515 => x"31544146",
   516 => x"20202036",
   517 => x"00000000",
   518 => x"20202e2e",
   519 => x"20202020",
   520 => x"00202020",
   521 => x"5c5b5e0e",
   522 => x"4a710e5d",
   523 => x"bfdce0c2",
   524 => x"7287cb02",
   525 => x"722bc74b",
   526 => x"9dffc14d",
   527 => x"4b7287c9",
   528 => x"4d722bc8",
   529 => x"c29dffc3",
   530 => x"83bfece4",
   531 => x"bfd4f2c0",
   532 => x"87d902ab",
   533 => x"5bd8f2c0",
   534 => x"1ed4d8c2",
   535 => x"caf04973",
   536 => x"7086c487",
   537 => x"87c50598",
   538 => x"e6c048c0",
   539 => x"dce0c287",
   540 => x"87d202bf",
   541 => x"91c44975",
   542 => x"81d4d8c2",
   543 => x"ffcf4c69",
   544 => x"9cffffff",
   545 => x"497587cb",
   546 => x"d8c291c2",
   547 => x"699f81d4",
   548 => x"2648744c",
   549 => x"264c264d",
   550 => x"0e4f264b",
   551 => x"5d5c5b5e",
   552 => x"cc86f40e",
   553 => x"66dc59a6",
   554 => x"dc87c702",
   555 => x"05bf9766",
   556 => x"48c087c5",
   557 => x"c887f4c2",
   558 => x"80c84866",
   559 => x"c0487e70",
   560 => x"49c11e78",
   561 => x"87d4c749",
   562 => x"4c7086c4",
   563 => x"fbc0029c",
   564 => x"e4e0c287",
   565 => x"4966dc4a",
   566 => x"87efdfff",
   567 => x"c0029870",
   568 => x"4a7487ea",
   569 => x"cb4966dc",
   570 => x"87d4e04b",
   571 => x"db029870",
   572 => x"741ec087",
   573 => x"87c4029c",
   574 => x"87c24dc0",
   575 => x"49754dc1",
   576 => x"c487d9c6",
   577 => x"9c4c7086",
   578 => x"87c5ff05",
   579 => x"c1029c74",
   580 => x"a4dc87d7",
   581 => x"69486e49",
   582 => x"49a4da78",
   583 => x"c44866c8",
   584 => x"58a6c880",
   585 => x"c448699f",
   586 => x"c2780866",
   587 => x"02bfdce0",
   588 => x"a4d487d2",
   589 => x"49699f49",
   590 => x"99ffffc0",
   591 => x"30d04871",
   592 => x"87c27e70",
   593 => x"486e7ec0",
   594 => x"80bf66c4",
   595 => x"780866c4",
   596 => x"c04866c8",
   597 => x"4966c878",
   598 => x"66c481cc",
   599 => x"66c879bf",
   600 => x"c081d049",
   601 => x"c248c179",
   602 => x"f448c087",
   603 => x"264d268e",
   604 => x"264b264c",
   605 => x"5b5e0e4f",
   606 => x"710e5d5c",
   607 => x"4d66d04c",
   608 => x"72496c4a",
   609 => x"c2b94da1",
   610 => x"4abfd8e0",
   611 => x"9972baff",
   612 => x"c0029971",
   613 => x"a4c487e4",
   614 => x"fa496b4b",
   615 => x"7b7087c6",
   616 => x"bfd4e0c2",
   617 => x"71816c49",
   618 => x"c2b9757c",
   619 => x"4abfd8e0",
   620 => x"9972baff",
   621 => x"ff059971",
   622 => x"7c7587dc",
   623 => x"4c264d26",
   624 => x"4f264b26",
   625 => x"711e731e",
   626 => x"f0e4c24b",
   627 => x"a3c449bf",
   628 => x"c24a6a4a",
   629 => x"d4e0c28a",
   630 => x"a17292bf",
   631 => x"d8e0c249",
   632 => x"9a6b4abf",
   633 => x"c049a172",
   634 => x"c859d8f2",
   635 => x"e9711e66",
   636 => x"86c487f9",
   637 => x"c4059870",
   638 => x"c248c087",
   639 => x"2648c187",
   640 => x"1e4f264b",
   641 => x"4b711e73",
   642 => x"e4c0029b",
   643 => x"c4e5c287",
   644 => x"c24a735b",
   645 => x"d4e0c28a",
   646 => x"c29249bf",
   647 => x"48bff0e4",
   648 => x"e5c28072",
   649 => x"487158c8",
   650 => x"e0c230c4",
   651 => x"edc058e4",
   652 => x"c0e5c287",
   653 => x"f4e4c248",
   654 => x"e5c278bf",
   655 => x"e4c248c4",
   656 => x"c278bff8",
   657 => x"02bfdce0",
   658 => x"e0c287c9",
   659 => x"c449bfd4",
   660 => x"c287c731",
   661 => x"49bffce4",
   662 => x"e0c231c4",
   663 => x"4b2659e4",
   664 => x"5e0e4f26",
   665 => x"710e5c5b",
   666 => x"724bc04a",
   667 => x"e0c0029a",
   668 => x"49a2da87",
   669 => x"c24b699f",
   670 => x"02bfdce0",
   671 => x"a2d487cf",
   672 => x"49699f49",
   673 => x"ffffc04c",
   674 => x"c234d09c",
   675 => x"744cc087",
   676 => x"fd4973b3",
   677 => x"4c2687ed",
   678 => x"4f264b26",
   679 => x"5c5b5e0e",
   680 => x"86f00e5d",
   681 => x"cf59a6c8",
   682 => x"f8ffffff",
   683 => x"c47ec04c",
   684 => x"87d80266",
   685 => x"48d0d8c2",
   686 => x"d8c278c0",
   687 => x"e5c248c8",
   688 => x"c278bfc4",
   689 => x"c248ccd8",
   690 => x"78bfc0e5",
   691 => x"48f1e0c2",
   692 => x"e0c250c0",
   693 => x"c249bfe0",
   694 => x"4abfd0d8",
   695 => x"c403aa71",
   696 => x"497287cb",
   697 => x"c00599cf",
   698 => x"f2c087e9",
   699 => x"d8c248d4",
   700 => x"c278bfc8",
   701 => x"c21ed4d8",
   702 => x"49bfc8d8",
   703 => x"48c8d8c2",
   704 => x"7178a1c1",
   705 => x"c487e4e5",
   706 => x"d0f2c086",
   707 => x"d4d8c248",
   708 => x"c087cc78",
   709 => x"48bfd0f2",
   710 => x"c080e0c0",
   711 => x"c258d4f2",
   712 => x"48bfd0d8",
   713 => x"d8c280c1",
   714 => x"902758d4",
   715 => x"bf00000c",
   716 => x"9d4dbf97",
   717 => x"87e5c202",
   718 => x"02ade5c3",
   719 => x"c087dec2",
   720 => x"4bbfd0f2",
   721 => x"1149a3cb",
   722 => x"05accf4c",
   723 => x"7587d2c1",
   724 => x"c199df49",
   725 => x"c291cd89",
   726 => x"c181e4e0",
   727 => x"51124aa3",
   728 => x"124aa3c3",
   729 => x"4aa3c551",
   730 => x"a3c75112",
   731 => x"c951124a",
   732 => x"51124aa3",
   733 => x"124aa3ce",
   734 => x"4aa3d051",
   735 => x"a3d25112",
   736 => x"d451124a",
   737 => x"51124aa3",
   738 => x"124aa3d6",
   739 => x"4aa3d851",
   740 => x"a3dc5112",
   741 => x"de51124a",
   742 => x"51124aa3",
   743 => x"fcc07ec1",
   744 => x"c8497487",
   745 => x"edc00599",
   746 => x"d0497487",
   747 => x"87d30599",
   748 => x"0266e0c0",
   749 => x"7387ccc0",
   750 => x"66e0c049",
   751 => x"0298700f",
   752 => x"6e87d3c0",
   753 => x"87c6c005",
   754 => x"48e4e0c2",
   755 => x"f2c050c0",
   756 => x"c248bfd0",
   757 => x"e0c287e9",
   758 => x"50c048f1",
   759 => x"e0e0c27e",
   760 => x"d8c249bf",
   761 => x"714abfd0",
   762 => x"f5fb04aa",
   763 => x"ffffcf87",
   764 => x"c24cf8ff",
   765 => x"05bfc4e5",
   766 => x"c287c8c0",
   767 => x"02bfdce0",
   768 => x"c287fac1",
   769 => x"49bfccd8",
   770 => x"c287d9f0",
   771 => x"c458d0d8",
   772 => x"d8c248a6",
   773 => x"c278bfcc",
   774 => x"02bfdce0",
   775 => x"c487dbc0",
   776 => x"99744966",
   777 => x"c002a974",
   778 => x"a6c887c8",
   779 => x"c078c048",
   780 => x"a6c887e7",
   781 => x"c078c148",
   782 => x"66c487df",
   783 => x"f8ffcf49",
   784 => x"c002a999",
   785 => x"a6cc87c8",
   786 => x"c078c048",
   787 => x"a6cc87c5",
   788 => x"c878c148",
   789 => x"66cc48a6",
   790 => x"0566c878",
   791 => x"c487dec0",
   792 => x"89c24966",
   793 => x"bfd4e0c2",
   794 => x"f0e4c291",
   795 => x"807148bf",
   796 => x"58ccd8c2",
   797 => x"48d0d8c2",
   798 => x"d5f978c0",
   799 => x"cf48c087",
   800 => x"f8ffffff",
   801 => x"268ef04c",
   802 => x"264c264d",
   803 => x"004f264b",
   804 => x"00000000",
   805 => x"ffffffff",
   806 => x"48d4ff1e",
   807 => x"6878ffc3",
   808 => x"1e4f2648",
   809 => x"c348d4ff",
   810 => x"d0ff78ff",
   811 => x"78e1c048",
   812 => x"d448d4ff",
   813 => x"1e4f2678",
   814 => x"c048d0ff",
   815 => x"4f2678e0",
   816 => x"87d4ff1e",
   817 => x"02994970",
   818 => x"fbc087c6",
   819 => x"87f105a9",
   820 => x"4f264871",
   821 => x"5c5b5e0e",
   822 => x"c04b710e",
   823 => x"87f8fe4c",
   824 => x"02994970",
   825 => x"c087f9c0",
   826 => x"c002a9ec",
   827 => x"fbc087f2",
   828 => x"ebc002a9",
   829 => x"b766cc87",
   830 => x"87c703ac",
   831 => x"c20266d0",
   832 => x"71537187",
   833 => x"87c20299",
   834 => x"cbfe84c1",
   835 => x"99497087",
   836 => x"c087cd02",
   837 => x"c702a9ec",
   838 => x"a9fbc087",
   839 => x"87d5ff05",
   840 => x"c30266d0",
   841 => x"7b97c087",
   842 => x"05a9ecc0",
   843 => x"4a7487c4",
   844 => x"4a7487c5",
   845 => x"728a0ac0",
   846 => x"264c2648",
   847 => x"1e4f264b",
   848 => x"7087d5fd",
   849 => x"f0c04a49",
   850 => x"87c904aa",
   851 => x"01aaf9c0",
   852 => x"f0c087c3",
   853 => x"aac1c18a",
   854 => x"c187c904",
   855 => x"c301aada",
   856 => x"8af7c087",
   857 => x"4f264872",
   858 => x"5c5b5e0e",
   859 => x"86f80e5d",
   860 => x"7ec04c71",
   861 => x"c087ecfc",
   862 => x"c8f8c04b",
   863 => x"c049bf97",
   864 => x"87cf04a9",
   865 => x"c187f9fc",
   866 => x"c8f8c083",
   867 => x"ab49bf97",
   868 => x"c087f106",
   869 => x"bf97c8f8",
   870 => x"fb87cf02",
   871 => x"497087fa",
   872 => x"87c60299",
   873 => x"05a9ecc0",
   874 => x"4bc087f1",
   875 => x"7087e9fb",
   876 => x"87e4fb4d",
   877 => x"fb58a6c8",
   878 => x"4a7087de",
   879 => x"a4c883c1",
   880 => x"49699749",
   881 => x"87da05ad",
   882 => x"9749a4c9",
   883 => x"66c44969",
   884 => x"87ce05a9",
   885 => x"9749a4ca",
   886 => x"05aa4969",
   887 => x"7ec187c4",
   888 => x"ecc087d0",
   889 => x"87c602ad",
   890 => x"05adfbc0",
   891 => x"4bc087c4",
   892 => x"026e7ec1",
   893 => x"fa87f5fe",
   894 => x"487387fd",
   895 => x"4d268ef8",
   896 => x"4b264c26",
   897 => x"00004f26",
   898 => x"1e731e00",
   899 => x"c84bd4ff",
   900 => x"d0ff4a66",
   901 => x"78c5c848",
   902 => x"c148d4ff",
   903 => x"7b1178d4",
   904 => x"f9058ac1",
   905 => x"48d0ff87",
   906 => x"4b2678c4",
   907 => x"5e0e4f26",
   908 => x"0e5d5c5b",
   909 => x"7e7186f8",
   910 => x"e5c21e6e",
   911 => x"dae949d4",
   912 => x"7086c487",
   913 => x"e4c40298",
   914 => x"c8e6c187",
   915 => x"496e4cbf",
   916 => x"c887d5fc",
   917 => x"987058a6",
   918 => x"c487c505",
   919 => x"78c148a6",
   920 => x"c548d0ff",
   921 => x"48d4ff78",
   922 => x"c478d5c1",
   923 => x"89c14966",
   924 => x"e6c131c6",
   925 => x"4abf97c0",
   926 => x"ffb07148",
   927 => x"ff7808d4",
   928 => x"78c448d0",
   929 => x"97d0e5c2",
   930 => x"99d049bf",
   931 => x"c587dd02",
   932 => x"48d4ff78",
   933 => x"c078d6c1",
   934 => x"48d4ff4a",
   935 => x"c178ffc3",
   936 => x"aae0c082",
   937 => x"ff87f204",
   938 => x"78c448d0",
   939 => x"c348d4ff",
   940 => x"d0ff78ff",
   941 => x"ff78c548",
   942 => x"d3c148d4",
   943 => x"ff78c178",
   944 => x"78c448d0",
   945 => x"06acb7c0",
   946 => x"c287cbc2",
   947 => x"4bbfdce5",
   948 => x"737e748c",
   949 => x"ddc1029b",
   950 => x"4dc0c887",
   951 => x"abb7c08b",
   952 => x"c887c603",
   953 => x"c04da3c0",
   954 => x"d0e5c24b",
   955 => x"d049bf97",
   956 => x"87cf0299",
   957 => x"e5c21ec0",
   958 => x"c7eb49d4",
   959 => x"7086c487",
   960 => x"c287d84c",
   961 => x"c21ed4d8",
   962 => x"ea49d4e5",
   963 => x"4c7087f6",
   964 => x"d8c21e75",
   965 => x"f0fb49d4",
   966 => x"7486c887",
   967 => x"87c5059c",
   968 => x"cac148c0",
   969 => x"c21ec187",
   970 => x"e949d4e5",
   971 => x"86c487c7",
   972 => x"fe059b73",
   973 => x"4c6e87e3",
   974 => x"06acb7c0",
   975 => x"e5c287d1",
   976 => x"78c048d4",
   977 => x"78c080d0",
   978 => x"e5c280f4",
   979 => x"c078bfe0",
   980 => x"fd01acb7",
   981 => x"d0ff87f5",
   982 => x"ff78c548",
   983 => x"d3c148d4",
   984 => x"ff78c078",
   985 => x"78c448d0",
   986 => x"c2c048c1",
   987 => x"f848c087",
   988 => x"264d268e",
   989 => x"264b264c",
   990 => x"5b5e0e4f",
   991 => x"fc0e5d5c",
   992 => x"c04d7186",
   993 => x"04ad4c4b",
   994 => x"c087e8c0",
   995 => x"741ee8f5",
   996 => x"87c4029c",
   997 => x"87c24ac0",
   998 => x"49724ac1",
   999 => x"c487fdeb",
  1000 => x"c17e7086",
  1001 => x"c2056e83",
  1002 => x"c14b7587",
  1003 => x"06ab7584",
  1004 => x"6e87d8ff",
  1005 => x"268efc48",
  1006 => x"264c264d",
  1007 => x"1e4f264b",
  1008 => x"66c44a71",
  1009 => x"7287c505",
  1010 => x"87e2f949",
  1011 => x"5e0e4f26",
  1012 => x"0e5d5c5b",
  1013 => x"4c7186fc",
  1014 => x"c291de49",
  1015 => x"714dc0e6",
  1016 => x"026d9785",
  1017 => x"c287dcc1",
  1018 => x"49bff0e5",
  1019 => x"fe718174",
  1020 => x"7e7087c7",
  1021 => x"c0029848",
  1022 => x"e5c287f2",
  1023 => x"4a704bf4",
  1024 => x"c4ff49cb",
  1025 => x"4b7487dd",
  1026 => x"e6c193cc",
  1027 => x"83c483cc",
  1028 => x"7bd0c1c1",
  1029 => x"c3c14974",
  1030 => x"7b7587fa",
  1031 => x"97c4e6c1",
  1032 => x"c21e49bf",
  1033 => x"fe49f4e5",
  1034 => x"86c487d5",
  1035 => x"c3c14974",
  1036 => x"49c087e2",
  1037 => x"87fdc4c1",
  1038 => x"48cce5c2",
  1039 => x"c04950c0",
  1040 => x"fc87e6e2",
  1041 => x"264d268e",
  1042 => x"264b264c",
  1043 => x"0000004f",
  1044 => x"64616f4c",
  1045 => x"2e676e69",
  1046 => x"00002e2e",
  1047 => x"61422080",
  1048 => x"00006b63",
  1049 => x"64616f4c",
  1050 => x"202e2a20",
  1051 => x"00000000",
  1052 => x"0000203a",
  1053 => x"61422080",
  1054 => x"00006b63",
  1055 => x"78452080",
  1056 => x"00007469",
  1057 => x"49204453",
  1058 => x"2e74696e",
  1059 => x"0000002e",
  1060 => x"00004b4f",
  1061 => x"544f4f42",
  1062 => x"20202020",
  1063 => x"004d4f52",
  1064 => x"711e731e",
  1065 => x"e5c2494b",
  1066 => x"7181bff0",
  1067 => x"7087cafb",
  1068 => x"c4029a4a",
  1069 => x"e9e64987",
  1070 => x"f0e5c287",
  1071 => x"7378c048",
  1072 => x"87fac149",
  1073 => x"4f264b26",
  1074 => x"711e731e",
  1075 => x"4aa3c44b",
  1076 => x"87d0c102",
  1077 => x"dc028ac1",
  1078 => x"c0028a87",
  1079 => x"058a87f2",
  1080 => x"c287d3c1",
  1081 => x"02bff0e5",
  1082 => x"4887cbc1",
  1083 => x"e5c288c1",
  1084 => x"c1c158f4",
  1085 => x"f0e5c287",
  1086 => x"89c649bf",
  1087 => x"59f4e5c2",
  1088 => x"03a9b7c0",
  1089 => x"c287efc0",
  1090 => x"c048f0e5",
  1091 => x"87e6c078",
  1092 => x"bfece5c2",
  1093 => x"c287df02",
  1094 => x"48bff0e5",
  1095 => x"e5c280c1",
  1096 => x"87d258f4",
  1097 => x"bfece5c2",
  1098 => x"c287cb02",
  1099 => x"48bff0e5",
  1100 => x"e5c280c6",
  1101 => x"497358f4",
  1102 => x"4b2687c4",
  1103 => x"5e0e4f26",
  1104 => x"0e5d5c5b",
  1105 => x"a6d086f0",
  1106 => x"d4d8c259",
  1107 => x"c24cc04d",
  1108 => x"c148ece5",
  1109 => x"48a6c878",
  1110 => x"7e7578c0",
  1111 => x"bff0e5c2",
  1112 => x"06a8c048",
  1113 => x"c887c0c1",
  1114 => x"7e755ca6",
  1115 => x"48d4d8c2",
  1116 => x"f2c00298",
  1117 => x"4d66c487",
  1118 => x"1ee8f5c0",
  1119 => x"c40266cc",
  1120 => x"c24cc087",
  1121 => x"744cc187",
  1122 => x"87d0e449",
  1123 => x"7e7086c4",
  1124 => x"66c885c1",
  1125 => x"cc80c148",
  1126 => x"e5c258a6",
  1127 => x"03adbff0",
  1128 => x"056e87c5",
  1129 => x"6e87d1ff",
  1130 => x"754cc04d",
  1131 => x"dcc3029d",
  1132 => x"e8f5c087",
  1133 => x"0266cc1e",
  1134 => x"a6c887c7",
  1135 => x"c578c048",
  1136 => x"48a6c887",
  1137 => x"66c878c1",
  1138 => x"87d0e349",
  1139 => x"7e7086c4",
  1140 => x"c2029848",
  1141 => x"cb4987e4",
  1142 => x"49699781",
  1143 => x"c10299d0",
  1144 => x"497487d4",
  1145 => x"e6c191cc",
  1146 => x"c2c181cc",
  1147 => x"81c879e0",
  1148 => x"7451ffc3",
  1149 => x"c291de49",
  1150 => x"714dc0e6",
  1151 => x"97c1c285",
  1152 => x"49a5c17d",
  1153 => x"c251e0c0",
  1154 => x"bf97e4e0",
  1155 => x"c187d202",
  1156 => x"4ba5c284",
  1157 => x"4ae4e0c2",
  1158 => x"fcfe49db",
  1159 => x"d9c187c5",
  1160 => x"49a5cd87",
  1161 => x"84c151c0",
  1162 => x"6e4ba5c2",
  1163 => x"fe49cb4a",
  1164 => x"c187f0fb",
  1165 => x"497487c4",
  1166 => x"e6c191cc",
  1167 => x"ffc081cc",
  1168 => x"e0c279ce",
  1169 => x"02bf97e4",
  1170 => x"497487d8",
  1171 => x"84c191de",
  1172 => x"4bc0e6c2",
  1173 => x"e0c28371",
  1174 => x"49dd4ae4",
  1175 => x"87c3fbfe",
  1176 => x"4b7487d8",
  1177 => x"e6c293de",
  1178 => x"a3cb83c0",
  1179 => x"c151c049",
  1180 => x"4a6e7384",
  1181 => x"fafe49cb",
  1182 => x"66c887e9",
  1183 => x"cc80c148",
  1184 => x"acc758a6",
  1185 => x"87c5c003",
  1186 => x"e4fc056e",
  1187 => x"03acc787",
  1188 => x"c287e4c0",
  1189 => x"c048ece5",
  1190 => x"cc497478",
  1191 => x"cce6c191",
  1192 => x"ceffc081",
  1193 => x"de497479",
  1194 => x"c0e6c291",
  1195 => x"c151c081",
  1196 => x"04acc784",
  1197 => x"c187dcff",
  1198 => x"c048e8e7",
  1199 => x"c180f750",
  1200 => x"c140e4cc",
  1201 => x"c878dcc1",
  1202 => x"c8c3c180",
  1203 => x"4966cc78",
  1204 => x"87c0f9c0",
  1205 => x"4d268ef0",
  1206 => x"4b264c26",
  1207 => x"731e4f26",
  1208 => x"494b711e",
  1209 => x"e6c191cc",
  1210 => x"a1c881cc",
  1211 => x"c0e6c14a",
  1212 => x"c9501248",
  1213 => x"f8c04aa1",
  1214 => x"501248c8",
  1215 => x"e6c181ca",
  1216 => x"501148c4",
  1217 => x"97c4e6c1",
  1218 => x"c01e49bf",
  1219 => x"87eff249",
  1220 => x"e9f84973",
  1221 => x"268efc87",
  1222 => x"1e4f264b",
  1223 => x"f9c049c0",
  1224 => x"4f2687d3",
  1225 => x"494a711e",
  1226 => x"e6c191cc",
  1227 => x"81c881cc",
  1228 => x"48cce5c2",
  1229 => x"f0c05011",
  1230 => x"f5fe49a2",
  1231 => x"49c087ce",
  1232 => x"2687e6d6",
  1233 => x"d4ff1e4f",
  1234 => x"7affc34a",
  1235 => x"c048d0ff",
  1236 => x"7ade78e1",
  1237 => x"c8487a71",
  1238 => x"7a7028b7",
  1239 => x"b7d04871",
  1240 => x"717a7028",
  1241 => x"28b7d848",
  1242 => x"d0ff7a70",
  1243 => x"78e0c048",
  1244 => x"5e0e4f26",
  1245 => x"0e5d5c5b",
  1246 => x"4d7186f4",
  1247 => x"c191cc49",
  1248 => x"c881cce6",
  1249 => x"a1ca4aa1",
  1250 => x"48a6c47e",
  1251 => x"bfc8e5c2",
  1252 => x"bf976e78",
  1253 => x"4c66c44b",
  1254 => x"48122c73",
  1255 => x"7058a6cc",
  1256 => x"c984c19c",
  1257 => x"49699781",
  1258 => x"c204acb7",
  1259 => x"6e4cc087",
  1260 => x"c84abf97",
  1261 => x"31724966",
  1262 => x"66c4b9ff",
  1263 => x"72487499",
  1264 => x"b14a7030",
  1265 => x"59cce5c2",
  1266 => x"87f9fd71",
  1267 => x"e5c21ec7",
  1268 => x"c11ebfe8",
  1269 => x"c21ecce6",
  1270 => x"bf97cce5",
  1271 => x"87f4c149",
  1272 => x"f4c04975",
  1273 => x"8ee887ee",
  1274 => x"4c264d26",
  1275 => x"4f264b26",
  1276 => x"711e731e",
  1277 => x"f9fd494b",
  1278 => x"fd497387",
  1279 => x"4b2687f4",
  1280 => x"731e4f26",
  1281 => x"c24b711e",
  1282 => x"d6024aa3",
  1283 => x"058ac187",
  1284 => x"c287e2c0",
  1285 => x"02bfe8e5",
  1286 => x"c14887db",
  1287 => x"ece5c288",
  1288 => x"c287d258",
  1289 => x"02bfece5",
  1290 => x"e5c287cb",
  1291 => x"c148bfe8",
  1292 => x"ece5c280",
  1293 => x"c21ec758",
  1294 => x"1ebfe8e5",
  1295 => x"1ecce6c1",
  1296 => x"97cce5c2",
  1297 => x"87cc49bf",
  1298 => x"f3c04973",
  1299 => x"8ef487c6",
  1300 => x"4f264b26",
  1301 => x"5c5b5e0e",
  1302 => x"ccff0e5d",
  1303 => x"a6e4c086",
  1304 => x"48a6cc59",
  1305 => x"80c478c0",
  1306 => x"80c478c0",
  1307 => x"7866c8c1",
  1308 => x"78c180c4",
  1309 => x"78c180c4",
  1310 => x"48ece5c2",
  1311 => x"e2e078c1",
  1312 => x"87fce087",
  1313 => x"7087d1e0",
  1314 => x"acfbc04c",
  1315 => x"87f3c102",
  1316 => x"0566e0c0",
  1317 => x"c187e8c1",
  1318 => x"c44a66c4",
  1319 => x"c17e6a82",
  1320 => x"6e48e4c1",
  1321 => x"20412049",
  1322 => x"c1511041",
  1323 => x"c14866c4",
  1324 => x"6a78decb",
  1325 => x"7481c749",
  1326 => x"66c4c151",
  1327 => x"c181c849",
  1328 => x"48a6d851",
  1329 => x"c4c178c2",
  1330 => x"81c94966",
  1331 => x"c4c151c0",
  1332 => x"81ca4966",
  1333 => x"1ec151c0",
  1334 => x"496a1ed8",
  1335 => x"dfff81c8",
  1336 => x"86c887f2",
  1337 => x"4866c8c1",
  1338 => x"c701a8c0",
  1339 => x"48a6d087",
  1340 => x"87cf78c1",
  1341 => x"4866c8c1",
  1342 => x"a6d888c1",
  1343 => x"ff87c458",
  1344 => x"7487fdde",
  1345 => x"dacd029c",
  1346 => x"4866d087",
  1347 => x"a866ccc1",
  1348 => x"87cfcd03",
  1349 => x"c048a6c8",
  1350 => x"ddff7e78",
  1351 => x"4c7087fa",
  1352 => x"05acd0c1",
  1353 => x"c487e7c2",
  1354 => x"786e48a6",
  1355 => x"7087d0e0",
  1356 => x"66cc487e",
  1357 => x"87c506a8",
  1358 => x"6e48a6cc",
  1359 => x"d7ddff78",
  1360 => x"c04c7087",
  1361 => x"c105acec",
  1362 => x"66d087ee",
  1363 => x"c191cc49",
  1364 => x"c48166c4",
  1365 => x"4d6a4aa1",
  1366 => x"6e4aa1c8",
  1367 => x"e4ccc152",
  1368 => x"f3dcff79",
  1369 => x"9c4c7087",
  1370 => x"c087d902",
  1371 => x"d302acfb",
  1372 => x"ff557487",
  1373 => x"7087e1dc",
  1374 => x"c7029c4c",
  1375 => x"acfbc087",
  1376 => x"87edff05",
  1377 => x"c255e0c0",
  1378 => x"97c055c1",
  1379 => x"66e0c07d",
  1380 => x"a866c448",
  1381 => x"d087db05",
  1382 => x"66d44866",
  1383 => x"87ca04a8",
  1384 => x"c14866d0",
  1385 => x"58a6d480",
  1386 => x"66d487c8",
  1387 => x"d888c148",
  1388 => x"dbff58a6",
  1389 => x"4c7087e2",
  1390 => x"05acd0c1",
  1391 => x"66dc87c9",
  1392 => x"c080c148",
  1393 => x"c158a6e0",
  1394 => x"fd02acd0",
  1395 => x"486e87d9",
  1396 => x"a866e0c0",
  1397 => x"87ebc905",
  1398 => x"48a6e4c0",
  1399 => x"487478c0",
  1400 => x"c888fbc0",
  1401 => x"987058a6",
  1402 => x"87ddc902",
  1403 => x"c888cb48",
  1404 => x"987058a6",
  1405 => x"87cfc102",
  1406 => x"c888c948",
  1407 => x"987058a6",
  1408 => x"87ffc302",
  1409 => x"c888c448",
  1410 => x"987058a6",
  1411 => x"4887cf02",
  1412 => x"a6c888c1",
  1413 => x"02987058",
  1414 => x"c887e8c3",
  1415 => x"a6c887dc",
  1416 => x"78f0c048",
  1417 => x"87f0d9ff",
  1418 => x"ecc04c70",
  1419 => x"c3c002ac",
  1420 => x"5ca6cc87",
  1421 => x"02acecc0",
  1422 => x"d9ff87cd",
  1423 => x"4c7087da",
  1424 => x"05acecc0",
  1425 => x"c087f3ff",
  1426 => x"c002acec",
  1427 => x"d9ff87c4",
  1428 => x"1ec087c6",
  1429 => x"66d81eca",
  1430 => x"c191cc49",
  1431 => x"714866cc",
  1432 => x"58a6cc80",
  1433 => x"c44866c8",
  1434 => x"58a6d080",
  1435 => x"49bf66cc",
  1436 => x"87e0d9ff",
  1437 => x"1ede1ec1",
  1438 => x"49bf66d4",
  1439 => x"87d4d9ff",
  1440 => x"497086d0",
  1441 => x"8808c048",
  1442 => x"58a6ecc0",
  1443 => x"c006a8c0",
  1444 => x"e8c087ee",
  1445 => x"a8dd4866",
  1446 => x"87e4c003",
  1447 => x"49bf66c4",
  1448 => x"8166e8c0",
  1449 => x"c051e0c0",
  1450 => x"c14966e8",
  1451 => x"bf66c481",
  1452 => x"51c1c281",
  1453 => x"4966e8c0",
  1454 => x"66c481c2",
  1455 => x"51c081bf",
  1456 => x"cbc1486e",
  1457 => x"496e78de",
  1458 => x"66d881c8",
  1459 => x"c9496e51",
  1460 => x"5166dc81",
  1461 => x"81ca496e",
  1462 => x"d85166c8",
  1463 => x"80c14866",
  1464 => x"d058a6dc",
  1465 => x"66d44866",
  1466 => x"cbc004a8",
  1467 => x"4866d087",
  1468 => x"a6d480c1",
  1469 => x"87d1c558",
  1470 => x"c14866d4",
  1471 => x"58a6d888",
  1472 => x"ff87c6c5",
  1473 => x"c087f8d8",
  1474 => x"ff58a6ec",
  1475 => x"c087f0d8",
  1476 => x"c058a6f0",
  1477 => x"c005a8ec",
  1478 => x"48a687c9",
  1479 => x"7866e8c0",
  1480 => x"ff87c4c0",
  1481 => x"d087f1d5",
  1482 => x"91cc4966",
  1483 => x"4866c4c1",
  1484 => x"a6c88071",
  1485 => x"4a66c458",
  1486 => x"66c482c8",
  1487 => x"c081ca49",
  1488 => x"c05166e8",
  1489 => x"c14966ec",
  1490 => x"66e8c081",
  1491 => x"7148c189",
  1492 => x"c1497030",
  1493 => x"7a977189",
  1494 => x"bfc8e5c2",
  1495 => x"66e8c049",
  1496 => x"4a6a9729",
  1497 => x"c0987148",
  1498 => x"c458a6f4",
  1499 => x"80c44866",
  1500 => x"c858a6cc",
  1501 => x"c04dbf66",
  1502 => x"6e4866e0",
  1503 => x"c5c002a8",
  1504 => x"c07ec087",
  1505 => x"7ec187c2",
  1506 => x"e0c01e6e",
  1507 => x"ff49751e",
  1508 => x"c887c1d5",
  1509 => x"c04c7086",
  1510 => x"c106acb7",
  1511 => x"857487d4",
  1512 => x"49bf66c8",
  1513 => x"7581e0c0",
  1514 => x"c1c14b89",
  1515 => x"fe714af0",
  1516 => x"c287f0e5",
  1517 => x"c07e7585",
  1518 => x"c14866e4",
  1519 => x"a6e8c080",
  1520 => x"66f0c058",
  1521 => x"7081c149",
  1522 => x"c5c002a9",
  1523 => x"c04dc087",
  1524 => x"4dc187c2",
  1525 => x"66cc1e75",
  1526 => x"e0c049bf",
  1527 => x"8966c481",
  1528 => x"66c81e71",
  1529 => x"ebd3ff49",
  1530 => x"c086c887",
  1531 => x"ff01a8b7",
  1532 => x"e4c087c5",
  1533 => x"d3c00266",
  1534 => x"4966c487",
  1535 => x"e4c081c9",
  1536 => x"66c45166",
  1537 => x"f2cdc148",
  1538 => x"87cec078",
  1539 => x"c94966c4",
  1540 => x"c451c281",
  1541 => x"cfc14866",
  1542 => x"66d078f0",
  1543 => x"a866d448",
  1544 => x"87cbc004",
  1545 => x"c14866d0",
  1546 => x"58a6d480",
  1547 => x"d487dac0",
  1548 => x"88c14866",
  1549 => x"c058a6d8",
  1550 => x"d2ff87cf",
  1551 => x"4c7087c2",
  1552 => x"ff87c6c0",
  1553 => x"7087f9d1",
  1554 => x"4866dc4c",
  1555 => x"e0c080c1",
  1556 => x"9c7458a6",
  1557 => x"87cbc002",
  1558 => x"c14866d0",
  1559 => x"04a866cc",
  1560 => x"d087f1f2",
  1561 => x"a8c74866",
  1562 => x"87e1c003",
  1563 => x"c24c66d0",
  1564 => x"c048ece5",
  1565 => x"cc497478",
  1566 => x"66c4c191",
  1567 => x"4aa1c481",
  1568 => x"52c04a6a",
  1569 => x"c784c179",
  1570 => x"e2ff04ac",
  1571 => x"66e0c087",
  1572 => x"87e2c002",
  1573 => x"4966c4c1",
  1574 => x"c181d4c1",
  1575 => x"c14a66c4",
  1576 => x"52c082dc",
  1577 => x"79e4ccc1",
  1578 => x"4966c4c1",
  1579 => x"c181d8c1",
  1580 => x"c079f4c1",
  1581 => x"c4c187d6",
  1582 => x"d4c14966",
  1583 => x"66c4c181",
  1584 => x"82d8c14a",
  1585 => x"7afcc1c1",
  1586 => x"79dbccc1",
  1587 => x"4966c4c1",
  1588 => x"c181e0c1",
  1589 => x"ff79c2d0",
  1590 => x"cc87dccf",
  1591 => x"ccff4866",
  1592 => x"264d268e",
  1593 => x"264b264c",
  1594 => x"1ec71e4f",
  1595 => x"bfe8e5c2",
  1596 => x"cce6c11e",
  1597 => x"cce5c21e",
  1598 => x"ed49bf97",
  1599 => x"e6c187d6",
  1600 => x"e1c049cc",
  1601 => x"8ef487dc",
  1602 => x"731e4f26",
  1603 => x"87d9c71e",
  1604 => x"48f4e5c2",
  1605 => x"d4ff50c0",
  1606 => x"78ffc348",
  1607 => x"49c4c2c1",
  1608 => x"87c3defe",
  1609 => x"87d8e9fe",
  1610 => x"cd029870",
  1611 => x"cbf1fe87",
  1612 => x"02987087",
  1613 => x"4ac187c4",
  1614 => x"4ac087c2",
  1615 => x"c8029a72",
  1616 => x"d0c2c187",
  1617 => x"deddfe49",
  1618 => x"e8e5c287",
  1619 => x"c278c048",
  1620 => x"c048cce5",
  1621 => x"d0fe4950",
  1622 => x"fcefc087",
  1623 => x"9b4b7087",
  1624 => x"c187cf02",
  1625 => x"c75be8e7",
  1626 => x"87e8de49",
  1627 => x"e0c049c1",
  1628 => x"eec287c3",
  1629 => x"e4e1c087",
  1630 => x"2687fa87",
  1631 => x"004f264b",
  1632 => x"00000000",
  1633 => x"00000000",
  1634 => x"00000001",
  1635 => x"00000fce",
  1636 => x"00002980",
  1637 => x"00000000",
  1638 => x"00000fce",
  1639 => x"0000299e",
  1640 => x"00000000",
  1641 => x"00000fce",
  1642 => x"000029bc",
  1643 => x"00000000",
  1644 => x"00000fce",
  1645 => x"000029da",
  1646 => x"00000000",
  1647 => x"00000fce",
  1648 => x"000029f8",
  1649 => x"00000000",
  1650 => x"00000fce",
  1651 => x"00002a16",
  1652 => x"00000000",
  1653 => x"00000fce",
  1654 => x"00002a34",
  1655 => x"00000000",
  1656 => x"00001324",
  1657 => x"00000000",
  1658 => x"00000000",
  1659 => x"000010c8",
  1660 => x"00000000",
  1661 => x"00000000",
  1662 => x"00001094",
  1663 => x"db86fc1e",
  1664 => x"fc7e7087",
  1665 => x"1e4f268e",
  1666 => x"c048f0fe",
  1667 => x"7909cd78",
  1668 => x"1e4f2609",
  1669 => x"49fce7c1",
  1670 => x"4f2687ed",
  1671 => x"bff0fe1e",
  1672 => x"1e4f2648",
  1673 => x"c148f0fe",
  1674 => x"1e4f2678",
  1675 => x"c048f0fe",
  1676 => x"1e4f2678",
  1677 => x"52c04a71",
  1678 => x"0e4f2651",
  1679 => x"5d5c5b5e",
  1680 => x"7186f40e",
  1681 => x"7e6d974d",
  1682 => x"974ca5c1",
  1683 => x"a6c8486c",
  1684 => x"c4486e58",
  1685 => x"c505a866",
  1686 => x"c048ff87",
  1687 => x"caff87e6",
  1688 => x"49a5c287",
  1689 => x"714b6c97",
  1690 => x"6b974ba3",
  1691 => x"7e6c974b",
  1692 => x"80c1486e",
  1693 => x"c758a6c8",
  1694 => x"58a6cc98",
  1695 => x"fe7c9770",
  1696 => x"487387e1",
  1697 => x"4d268ef4",
  1698 => x"4b264c26",
  1699 => x"5e0e4f26",
  1700 => x"f40e5c5b",
  1701 => x"d84c7186",
  1702 => x"ffc34a66",
  1703 => x"4ba4c29a",
  1704 => x"73496c97",
  1705 => x"517249a1",
  1706 => x"6e7e6c97",
  1707 => x"c880c148",
  1708 => x"98c758a6",
  1709 => x"7058a6cc",
  1710 => x"268ef454",
  1711 => x"264b264c",
  1712 => x"86fc1e4f",
  1713 => x"e087e4fd",
  1714 => x"c0494abf",
  1715 => x"0299c0e0",
  1716 => x"1e7287cb",
  1717 => x"49e8e9c2",
  1718 => x"c487f3fe",
  1719 => x"87fcfc86",
  1720 => x"fefc7e70",
  1721 => x"268efc87",
  1722 => x"e9c21e4f",
  1723 => x"c2fd49e8",
  1724 => x"c1ebc187",
  1725 => x"87cffc49",
  1726 => x"2687edc4",
  1727 => x"5b5e0e4f",
  1728 => x"fc0e5d5c",
  1729 => x"ff7e7186",
  1730 => x"e9c24dd4",
  1731 => x"eafc49e8",
  1732 => x"c04b7087",
  1733 => x"c204abb7",
  1734 => x"f0c387f8",
  1735 => x"87c905ab",
  1736 => x"48e0efc1",
  1737 => x"d9c278c1",
  1738 => x"abe0c387",
  1739 => x"c187c905",
  1740 => x"c148e4ef",
  1741 => x"87cac278",
  1742 => x"bfe4efc1",
  1743 => x"c287c602",
  1744 => x"c24ca3c0",
  1745 => x"c14c7387",
  1746 => x"02bfe0ef",
  1747 => x"7487e0c0",
  1748 => x"29b7c449",
  1749 => x"e8efc191",
  1750 => x"cf4a7481",
  1751 => x"c192c29a",
  1752 => x"70307248",
  1753 => x"72baff4a",
  1754 => x"70986948",
  1755 => x"7487db79",
  1756 => x"29b7c449",
  1757 => x"e8efc191",
  1758 => x"cf4a7481",
  1759 => x"c392c29a",
  1760 => x"70307248",
  1761 => x"b069484a",
  1762 => x"056e7970",
  1763 => x"ff87e7c0",
  1764 => x"e1c848d0",
  1765 => x"c17dc578",
  1766 => x"02bfe4ef",
  1767 => x"e0c387c3",
  1768 => x"e0efc17d",
  1769 => x"87c302bf",
  1770 => x"737df0c3",
  1771 => x"48d0ff7d",
  1772 => x"c078e1c8",
  1773 => x"efc178e0",
  1774 => x"78c048e4",
  1775 => x"48e0efc1",
  1776 => x"e9c278c0",
  1777 => x"f2f949e8",
  1778 => x"c04b7087",
  1779 => x"fd03abb7",
  1780 => x"48c087c8",
  1781 => x"4d268efc",
  1782 => x"4b264c26",
  1783 => x"00004f26",
  1784 => x"00000000",
  1785 => x"00000000",
  1786 => x"00000000",
  1787 => x"00000000",
  1788 => x"00000000",
  1789 => x"00000000",
  1790 => x"00000000",
  1791 => x"00000000",
  1792 => x"00000000",
  1793 => x"00000000",
  1794 => x"00000000",
  1795 => x"00000000",
  1796 => x"00000000",
  1797 => x"00000000",
  1798 => x"00000000",
  1799 => x"00000000",
  1800 => x"00000000",
  1801 => x"00000000",
  1802 => x"724ac01e",
  1803 => x"c191c449",
  1804 => x"c081e8ef",
  1805 => x"d082c179",
  1806 => x"ee04aab7",
  1807 => x"0e4f2687",
  1808 => x"5d5c5b5e",
  1809 => x"f74d710e",
  1810 => x"4a7587e1",
  1811 => x"922ab7c4",
  1812 => x"82e8efc1",
  1813 => x"9ccf4c75",
  1814 => x"496a94c2",
  1815 => x"c32b744b",
  1816 => x"7448c29b",
  1817 => x"ff4c7030",
  1818 => x"714874bc",
  1819 => x"f67a7098",
  1820 => x"487387f1",
  1821 => x"4c264d26",
  1822 => x"4f264b26",
  1823 => x"48d0ff1e",
  1824 => x"7178e1c8",
  1825 => x"08d4ff48",
  1826 => x"4866c478",
  1827 => x"7808d4ff",
  1828 => x"711e4f26",
  1829 => x"4966c44a",
  1830 => x"ff49721e",
  1831 => x"d0ff87de",
  1832 => x"78e0c048",
  1833 => x"4f268efc",
  1834 => x"711e731e",
  1835 => x"4966c84b",
  1836 => x"c14a731e",
  1837 => x"ff49a2e0",
  1838 => x"8efc87d8",
  1839 => x"4f264b26",
  1840 => x"48d0ff1e",
  1841 => x"7178c9c8",
  1842 => x"08d4ff48",
  1843 => x"1e4f2678",
  1844 => x"eb494a71",
  1845 => x"48d0ff87",
  1846 => x"4f2678c8",
  1847 => x"711e731e",
  1848 => x"c0eac24b",
  1849 => x"87c302bf",
  1850 => x"ff87ebc2",
  1851 => x"c9c848d0",
  1852 => x"c0487378",
  1853 => x"d4ffb0e0",
  1854 => x"e9c27808",
  1855 => x"78c048f4",
  1856 => x"c50266c8",
  1857 => x"49ffc387",
  1858 => x"49c087c2",
  1859 => x"59fce9c2",
  1860 => x"c60266cc",
  1861 => x"d5d5c587",
  1862 => x"cf87c44a",
  1863 => x"c24affff",
  1864 => x"c25ac0ea",
  1865 => x"c148c0ea",
  1866 => x"264b2678",
  1867 => x"5b5e0e4f",
  1868 => x"710e5d5c",
  1869 => x"fce9c24d",
  1870 => x"9d754bbf",
  1871 => x"4987cb02",
  1872 => x"f3c191c8",
  1873 => x"82714ad4",
  1874 => x"f7c187c4",
  1875 => x"4cc04ad4",
  1876 => x"99734912",
  1877 => x"bff8e9c2",
  1878 => x"ffb87148",
  1879 => x"c17808d4",
  1880 => x"c8842bb7",
  1881 => x"e704acb7",
  1882 => x"f4e9c287",
  1883 => x"80c848bf",
  1884 => x"58f8e9c2",
  1885 => x"4c264d26",
  1886 => x"4f264b26",
  1887 => x"711e731e",
  1888 => x"9a4a134b",
  1889 => x"7287cb02",
  1890 => x"87e1fe49",
  1891 => x"059a4a13",
  1892 => x"4b2687f5",
  1893 => x"c21e4f26",
  1894 => x"49bff4e9",
  1895 => x"48f4e9c2",
  1896 => x"c478a1c1",
  1897 => x"03a9b7c0",
  1898 => x"d4ff87db",
  1899 => x"f8e9c248",
  1900 => x"e9c278bf",
  1901 => x"c249bff4",
  1902 => x"c148f4e9",
  1903 => x"c0c478a1",
  1904 => x"e504a9b7",
  1905 => x"48d0ff87",
  1906 => x"eac278c8",
  1907 => x"78c048c0",
  1908 => x"00004f26",
  1909 => x"00000000",
  1910 => x"00000000",
  1911 => x"5f000000",
  1912 => x"0000005f",
  1913 => x"00030300",
  1914 => x"00000303",
  1915 => x"147f7f14",
  1916 => x"00147f7f",
  1917 => x"6b2e2400",
  1918 => x"00123a6b",
  1919 => x"18366a4c",
  1920 => x"0032566c",
  1921 => x"594f7e30",
  1922 => x"40683a77",
  1923 => x"07040000",
  1924 => x"00000003",
  1925 => x"3e1c0000",
  1926 => x"00004163",
  1927 => x"63410000",
  1928 => x"00001c3e",
  1929 => x"1c3e2a08",
  1930 => x"082a3e1c",
  1931 => x"3e080800",
  1932 => x"0008083e",
  1933 => x"e0800000",
  1934 => x"00000060",
  1935 => x"08080800",
  1936 => x"00080808",
  1937 => x"60000000",
  1938 => x"00000060",
  1939 => x"18306040",
  1940 => x"0103060c",
  1941 => x"597f3e00",
  1942 => x"003e7f4d",
  1943 => x"7f060400",
  1944 => x"0000007f",
  1945 => x"71634200",
  1946 => x"00464f59",
  1947 => x"49632200",
  1948 => x"00367f49",
  1949 => x"13161c18",
  1950 => x"00107f7f",
  1951 => x"45672700",
  1952 => x"00397d45",
  1953 => x"4b7e3c00",
  1954 => x"00307949",
  1955 => x"71010100",
  1956 => x"00070f79",
  1957 => x"497f3600",
  1958 => x"00367f49",
  1959 => x"494f0600",
  1960 => x"001e3f69",
  1961 => x"66000000",
  1962 => x"00000066",
  1963 => x"e6800000",
  1964 => x"00000066",
  1965 => x"14080800",
  1966 => x"00222214",
  1967 => x"14141400",
  1968 => x"00141414",
  1969 => x"14222200",
  1970 => x"00080814",
  1971 => x"51030200",
  1972 => x"00060f59",
  1973 => x"5d417f3e",
  1974 => x"001e1f55",
  1975 => x"097f7e00",
  1976 => x"007e7f09",
  1977 => x"497f7f00",
  1978 => x"00367f49",
  1979 => x"633e1c00",
  1980 => x"00414141",
  1981 => x"417f7f00",
  1982 => x"001c3e63",
  1983 => x"497f7f00",
  1984 => x"00414149",
  1985 => x"097f7f00",
  1986 => x"00010109",
  1987 => x"417f3e00",
  1988 => x"007a7b49",
  1989 => x"087f7f00",
  1990 => x"007f7f08",
  1991 => x"7f410000",
  1992 => x"0000417f",
  1993 => x"40602000",
  1994 => x"003f7f40",
  1995 => x"1c087f7f",
  1996 => x"00416336",
  1997 => x"407f7f00",
  1998 => x"00404040",
  1999 => x"0c067f7f",
  2000 => x"007f7f06",
  2001 => x"0c067f7f",
  2002 => x"007f7f18",
  2003 => x"417f3e00",
  2004 => x"003e7f41",
  2005 => x"097f7f00",
  2006 => x"00060f09",
  2007 => x"61417f3e",
  2008 => x"00407e7f",
  2009 => x"097f7f00",
  2010 => x"00667f19",
  2011 => x"4d6f2600",
  2012 => x"00327b59",
  2013 => x"7f010100",
  2014 => x"0001017f",
  2015 => x"407f3f00",
  2016 => x"003f7f40",
  2017 => x"703f0f00",
  2018 => x"000f3f70",
  2019 => x"18307f7f",
  2020 => x"007f7f30",
  2021 => x"1c366341",
  2022 => x"4163361c",
  2023 => x"7c060301",
  2024 => x"0103067c",
  2025 => x"4d597161",
  2026 => x"00414347",
  2027 => x"7f7f0000",
  2028 => x"00004141",
  2029 => x"0c060301",
  2030 => x"40603018",
  2031 => x"41410000",
  2032 => x"00007f7f",
  2033 => x"03060c08",
  2034 => x"00080c06",
  2035 => x"80808080",
  2036 => x"00808080",
  2037 => x"03000000",
  2038 => x"00000407",
  2039 => x"54742000",
  2040 => x"00787c54",
  2041 => x"447f7f00",
  2042 => x"00387c44",
  2043 => x"447c3800",
  2044 => x"00004444",
  2045 => x"447c3800",
  2046 => x"007f7f44",
  2047 => x"547c3800",
  2048 => x"00185c54",
  2049 => x"7f7e0400",
  2050 => x"00000505",
  2051 => x"a4bc1800",
  2052 => x"007cfca4",
  2053 => x"047f7f00",
  2054 => x"00787c04",
  2055 => x"3d000000",
  2056 => x"0000407d",
  2057 => x"80808000",
  2058 => x"00007dfd",
  2059 => x"107f7f00",
  2060 => x"00446c38",
  2061 => x"3f000000",
  2062 => x"0000407f",
  2063 => x"180c7c7c",
  2064 => x"00787c0c",
  2065 => x"047c7c00",
  2066 => x"00787c04",
  2067 => x"447c3800",
  2068 => x"00387c44",
  2069 => x"24fcfc00",
  2070 => x"00183c24",
  2071 => x"243c1800",
  2072 => x"00fcfc24",
  2073 => x"047c7c00",
  2074 => x"00080c04",
  2075 => x"545c4800",
  2076 => x"00207454",
  2077 => x"7f3f0400",
  2078 => x"00004444",
  2079 => x"407c3c00",
  2080 => x"007c7c40",
  2081 => x"603c1c00",
  2082 => x"001c3c60",
  2083 => x"30607c3c",
  2084 => x"003c7c60",
  2085 => x"10386c44",
  2086 => x"00446c38",
  2087 => x"e0bc1c00",
  2088 => x"001c3c60",
  2089 => x"74644400",
  2090 => x"00444c5c",
  2091 => x"3e080800",
  2092 => x"00414177",
  2093 => x"7f000000",
  2094 => x"0000007f",
  2095 => x"77414100",
  2096 => x"0008083e",
  2097 => x"03010102",
  2098 => x"00010202",
  2099 => x"7f7f7f7f",
  2100 => x"007f7f7f",
  2101 => x"1c1c0808",
  2102 => x"7f7f3e3e",
  2103 => x"3e3e7f7f",
  2104 => x"08081c1c",
  2105 => x"7c181000",
  2106 => x"0010187c",
  2107 => x"7c301000",
  2108 => x"0010307c",
  2109 => x"60603010",
  2110 => x"00061e78",
  2111 => x"183c6642",
  2112 => x"0042663c",
  2113 => x"c26a3878",
  2114 => x"00386cc6",
  2115 => x"60000060",
  2116 => x"00600000",
  2117 => x"5c5b5e0e",
  2118 => x"86fc0e5d",
  2119 => x"eac27e71",
  2120 => x"c04cbfc8",
  2121 => x"c41ec04b",
  2122 => x"c402ab66",
  2123 => x"c24dc087",
  2124 => x"754dc187",
  2125 => x"ee49731e",
  2126 => x"86c887e2",
  2127 => x"ef49e0c0",
  2128 => x"a4c487eb",
  2129 => x"f0496a4a",
  2130 => x"c9f187f2",
  2131 => x"c184cc87",
  2132 => x"abb7c883",
  2133 => x"87cdff04",
  2134 => x"4d268efc",
  2135 => x"4b264c26",
  2136 => x"711e4f26",
  2137 => x"cceac24a",
  2138 => x"cceac25a",
  2139 => x"4978c748",
  2140 => x"2687e1fe",
  2141 => x"1e731e4f",
  2142 => x"b7c04a71",
  2143 => x"87d303aa",
  2144 => x"bff0d4c2",
  2145 => x"c187c405",
  2146 => x"c087c24b",
  2147 => x"f4d4c24b",
  2148 => x"c287c45b",
  2149 => x"fc5af4d4",
  2150 => x"f0d4c248",
  2151 => x"c14a78bf",
  2152 => x"a2c0c19a",
  2153 => x"87e7ec49",
  2154 => x"4f264b26",
  2155 => x"c44a711e",
  2156 => x"49721e66",
  2157 => x"fc87f1eb",
  2158 => x"1e4f268e",
  2159 => x"c348d4ff",
  2160 => x"d0ff78ff",
  2161 => x"78e1c048",
  2162 => x"c148d4ff",
  2163 => x"c4487178",
  2164 => x"08d4ff30",
  2165 => x"48d0ff78",
  2166 => x"2678e0c0",
  2167 => x"5b5e0e4f",
  2168 => x"f00e5d5c",
  2169 => x"48a6c886",
  2170 => x"bfec78c0",
  2171 => x"c280fc7e",
  2172 => x"78bfc8ea",
  2173 => x"bfd0eac2",
  2174 => x"4cbfe84d",
  2175 => x"bff0d4c2",
  2176 => x"87f9e349",
  2177 => x"f6e849c7",
  2178 => x"c2497087",
  2179 => x"87cf0599",
  2180 => x"bfe8d4c2",
  2181 => x"6eb9ff49",
  2182 => x"0299c199",
  2183 => x"cb87c0c2",
  2184 => x"cfcc49ee",
  2185 => x"58a6d087",
  2186 => x"d2e849c7",
  2187 => x"05987087",
  2188 => x"496e87c8",
  2189 => x"c10299c1",
  2190 => x"66cc87c2",
  2191 => x"7ebfec4b",
  2192 => x"bff0d4c2",
  2193 => x"87f5e249",
  2194 => x"f3cb4973",
  2195 => x"02987087",
  2196 => x"d4c287d7",
  2197 => x"c149bfd0",
  2198 => x"d4d4c2b9",
  2199 => x"dafd7159",
  2200 => x"49eecb87",
  2201 => x"7087cdcb",
  2202 => x"e749c74b",
  2203 => x"987087d1",
  2204 => x"87c9ff05",
  2205 => x"99c1496e",
  2206 => x"87c1ff05",
  2207 => x"bff0d4c2",
  2208 => x"c2bac14a",
  2209 => x"fc5af4d4",
  2210 => x"c10a7a0a",
  2211 => x"a2c0c19a",
  2212 => x"87fbe849",
  2213 => x"e649dac1",
  2214 => x"a6c887e5",
  2215 => x"c278c148",
  2216 => x"6e48e8d4",
  2217 => x"f0d4c278",
  2218 => x"c7c105bf",
  2219 => x"c0c0c887",
  2220 => x"c8d7c24b",
  2221 => x"49154d7e",
  2222 => x"87c3e649",
  2223 => x"c0029870",
  2224 => x"b47387c2",
  2225 => x"052bb7c1",
  2226 => x"7487ebff",
  2227 => x"99ffc349",
  2228 => x"49c01e71",
  2229 => x"7487d5fb",
  2230 => x"29b7c849",
  2231 => x"49c11e71",
  2232 => x"c887c9fb",
  2233 => x"49fdc386",
  2234 => x"c387d4e5",
  2235 => x"cee549fa",
  2236 => x"87d1c887",
  2237 => x"ffc34974",
  2238 => x"2cb7c899",
  2239 => x"9c74b471",
  2240 => x"ff87df02",
  2241 => x"497ebfc8",
  2242 => x"bfecd4c2",
  2243 => x"a9e0c289",
  2244 => x"87c5c003",
  2245 => x"cfc04cc0",
  2246 => x"ecd4c287",
  2247 => x"c0786e48",
  2248 => x"d4c287c6",
  2249 => x"78c048ec",
  2250 => x"99c84974",
  2251 => x"87cec005",
  2252 => x"e449f5c3",
  2253 => x"497087c9",
  2254 => x"c00299c2",
  2255 => x"eac287ea",
  2256 => x"c002bfcc",
  2257 => x"c14887ca",
  2258 => x"d0eac288",
  2259 => x"87d3c058",
  2260 => x"c14866c4",
  2261 => x"7e7080e0",
  2262 => x"c002bf6e",
  2263 => x"ff4b87c5",
  2264 => x"c80f7349",
  2265 => x"78c148a6",
  2266 => x"99c44974",
  2267 => x"87cec005",
  2268 => x"e349f2c3",
  2269 => x"497087c9",
  2270 => x"c00299c2",
  2271 => x"eac287f0",
  2272 => x"487ebfcc",
  2273 => x"03a8b7c7",
  2274 => x"6e87cbc0",
  2275 => x"c280c148",
  2276 => x"c058d0ea",
  2277 => x"66c487d3",
  2278 => x"80e0c148",
  2279 => x"bf6e7e70",
  2280 => x"87c5c002",
  2281 => x"7349fe4b",
  2282 => x"48a6c80f",
  2283 => x"fdc378c1",
  2284 => x"87cbe249",
  2285 => x"99c24970",
  2286 => x"87e6c002",
  2287 => x"bfcceac2",
  2288 => x"87c9c002",
  2289 => x"48cceac2",
  2290 => x"d0c078c0",
  2291 => x"4a66c487",
  2292 => x"6a82e0c1",
  2293 => x"87c5c002",
  2294 => x"7349fd4b",
  2295 => x"48a6c80f",
  2296 => x"fac378c1",
  2297 => x"87d7e149",
  2298 => x"99c24970",
  2299 => x"87edc002",
  2300 => x"bfcceac2",
  2301 => x"a8b7c748",
  2302 => x"87c9c003",
  2303 => x"48cceac2",
  2304 => x"d3c078c7",
  2305 => x"4866c487",
  2306 => x"7080e0c1",
  2307 => x"02bf6e7e",
  2308 => x"4b87c5c0",
  2309 => x"0f7349fc",
  2310 => x"c148a6c8",
  2311 => x"c3487478",
  2312 => x"7e7098f0",
  2313 => x"c0059848",
  2314 => x"dac187ce",
  2315 => x"87cfe049",
  2316 => x"99c24970",
  2317 => x"87d0c202",
  2318 => x"c349eecb",
  2319 => x"a6d087f6",
  2320 => x"c4eac258",
  2321 => x"c250c048",
  2322 => x"bf97c4ea",
  2323 => x"87d8c105",
  2324 => x"cdc0056e",
  2325 => x"49dac187",
  2326 => x"87e3dfff",
  2327 => x"c1029870",
  2328 => x"bfe887c6",
  2329 => x"ffc3494b",
  2330 => x"2bb7c899",
  2331 => x"d4c2b371",
  2332 => x"ff49bff0",
  2333 => x"cc87c6da",
  2334 => x"c3c34966",
  2335 => x"02987087",
  2336 => x"c287c6c0",
  2337 => x"c148c4ea",
  2338 => x"c4eac250",
  2339 => x"c005bf97",
  2340 => x"497387d6",
  2341 => x"0599f0c3",
  2342 => x"c187c7ff",
  2343 => x"deff49da",
  2344 => x"987087dd",
  2345 => x"87fafe05",
  2346 => x"c248a6cc",
  2347 => x"78bfccea",
  2348 => x"cc4966cc",
  2349 => x"4866c491",
  2350 => x"7e708071",
  2351 => x"c002bf6e",
  2352 => x"cc4b87c6",
  2353 => x"0f734966",
  2354 => x"c0029d75",
  2355 => x"026d87e9",
  2356 => x"6d87e4c0",
  2357 => x"e6ddff49",
  2358 => x"c1497087",
  2359 => x"cbc00299",
  2360 => x"4ba5c487",
  2361 => x"bfcceac2",
  2362 => x"0f4b6b49",
  2363 => x"c00285c8",
  2364 => x"056d87c5",
  2365 => x"c887dcff",
  2366 => x"c8c00266",
  2367 => x"cceac287",
  2368 => x"cff049bf",
  2369 => x"268ef087",
  2370 => x"264c264d",
  2371 => x"004f264b",
  2372 => x"00000000",
  2373 => x"00000010",
  2374 => x"14111258",
  2375 => x"231c1b1d",
  2376 => x"9491595a",
  2377 => x"f4ebf2f5",
  2378 => x"00000000",
  2379 => x"00000000",
  2380 => x"00000000",
  2381 => x"ff4a711e",
  2382 => x"7249bfc8",
  2383 => x"4f2648a1",
  2384 => x"bfc8ff1e",
  2385 => x"c0c0fe89",
  2386 => x"a9c0c0c0",
  2387 => x"c087c401",
  2388 => x"c187c24a",
  2389 => x"2648724a",
  2390 => x"1e731e4f",
  2391 => x"e6c14bc0",
  2392 => x"50c048c0",
  2393 => x"bfd8d7c2",
  2394 => x"c1e3fe49",
  2395 => x"05987087",
  2396 => x"d6c287c4",
  2397 => x"e6c14bcc",
  2398 => x"50c148c0",
  2399 => x"bfdcd7c2",
  2400 => x"e9e2fe49",
  2401 => x"26487387",
  2402 => x"004f264b",
  2403 => x"5f434247",
  2404 => x"534f4942",
  2405 => x"4e49422e",
  2406 => x"746f6e20",
  2407 => x"756f6620",
  2408 => x"6f20646e",
  2409 => x"4453206e",
  2410 => x"72616320",
  2411 => x"00000064",
  2412 => x"5f434247",
  2413 => x"534f4942",
  2414 => x"004e4942",
  2415 => x"4f545541",
  2416 => x"544f4f42",
  2417 => x"00004247",
  2418 => x"11141258",
  2419 => x"231c1b1d",
  2420 => x"9194595a",
  2421 => x"f4ebf2f5",
  2422 => x"000025b0",
  2423 => x"000025bc",
  2424 => x"00001a13",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
