
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"f4",x"e8",x"c2",x"87"),
    12 => (x"48",x"c0",x"c8",x"4e"),
    13 => (x"d5",x"c1",x"28",x"c2"),
    14 => (x"ea",x"d6",x"e5",x"ea"),
    15 => (x"c1",x"46",x"71",x"49"),
    16 => (x"87",x"f9",x"01",x"88"),
    17 => (x"49",x"f4",x"e8",x"c2"),
    18 => (x"48",x"c4",x"d6",x"c2"),
    19 => (x"03",x"89",x"d0",x"89"),
    20 => (x"40",x"40",x"40",x"c0"),
    21 => (x"d0",x"87",x"f6",x"40"),
    22 => (x"50",x"c0",x"05",x"81"),
    23 => (x"f9",x"05",x"89",x"c1"),
    24 => (x"c3",x"d6",x"c2",x"87"),
    25 => (x"ff",x"d5",x"c2",x"4d"),
    26 => (x"02",x"ad",x"74",x"4c"),
    27 => (x"0f",x"24",x"87",x"c4"),
    28 => (x"e2",x"c1",x"87",x"f7"),
    29 => (x"d6",x"c2",x"87",x"d8"),
    30 => (x"d6",x"c2",x"4d",x"c3"),
    31 => (x"ad",x"74",x"4c",x"c3"),
    32 => (x"c4",x"87",x"c6",x"02"),
    33 => (x"f5",x"0f",x"6c",x"8c"),
    34 => (x"87",x"fd",x"00",x"87"),
    35 => (x"71",x"86",x"fc",x"1e"),
    36 => (x"49",x"c0",x"ff",x"4a"),
    37 => (x"c0",x"c4",x"48",x"69"),
    38 => (x"48",x"7e",x"70",x"98"),
    39 => (x"87",x"f4",x"02",x"98"),
    40 => (x"fc",x"48",x"79",x"72"),
    41 => (x"0e",x"4f",x"26",x"8e"),
    42 => (x"0e",x"5c",x"5b",x"5e"),
    43 => (x"4c",x"c0",x"4b",x"71"),
    44 => (x"02",x"9a",x"4a",x"13"),
    45 => (x"49",x"72",x"87",x"cd"),
    46 => (x"c1",x"87",x"d1",x"ff"),
    47 => (x"9a",x"4a",x"13",x"84"),
    48 => (x"74",x"87",x"f3",x"05"),
    49 => (x"26",x"4c",x"26",x"48"),
    50 => (x"1e",x"4f",x"26",x"4b"),
    51 => (x"1e",x"73",x"1e",x"72"),
    52 => (x"02",x"11",x"48",x"12"),
    53 => (x"c3",x"4b",x"87",x"ca"),
    54 => (x"73",x"9b",x"98",x"df"),
    55 => (x"87",x"f0",x"02",x"88"),
    56 => (x"4a",x"26",x"4b",x"26"),
    57 => (x"73",x"1e",x"4f",x"26"),
    58 => (x"c1",x"1e",x"72",x"1e"),
    59 => (x"87",x"ca",x"04",x"8b"),
    60 => (x"02",x"11",x"48",x"12"),
    61 => (x"02",x"88",x"87",x"c4"),
    62 => (x"4a",x"26",x"87",x"f1"),
    63 => (x"4f",x"26",x"4b",x"26"),
    64 => (x"73",x"1e",x"74",x"1e"),
    65 => (x"c1",x"1e",x"72",x"1e"),
    66 => (x"87",x"cf",x"04",x"8b"),
    67 => (x"02",x"11",x"48",x"12"),
    68 => (x"df",x"4c",x"87",x"c9"),
    69 => (x"88",x"74",x"9c",x"98"),
    70 => (x"26",x"87",x"ec",x"02"),
    71 => (x"26",x"4b",x"26",x"4a"),
    72 => (x"1e",x"4f",x"26",x"4c"),
    73 => (x"73",x"81",x"48",x"73"),
    74 => (x"87",x"c5",x"02",x"a9"),
    75 => (x"f6",x"05",x"53",x"12"),
    76 => (x"0e",x"4f",x"26",x"87"),
    77 => (x"0e",x"5c",x"5b",x"5e"),
    78 => (x"d4",x"ff",x"4a",x"71"),
    79 => (x"4b",x"66",x"cc",x"4c"),
    80 => (x"71",x"8b",x"c1",x"49"),
    81 => (x"87",x"ce",x"02",x"99"),
    82 => (x"6c",x"7c",x"ff",x"c3"),
    83 => (x"c1",x"49",x"73",x"52"),
    84 => (x"05",x"99",x"71",x"8b"),
    85 => (x"4c",x"26",x"87",x"f2"),
    86 => (x"4f",x"26",x"4b",x"26"),
    87 => (x"ff",x"1e",x"73",x"1e"),
    88 => (x"ff",x"c3",x"4b",x"d4"),
    89 => (x"c3",x"4a",x"6b",x"7b"),
    90 => (x"49",x"6b",x"7b",x"ff"),
    91 => (x"b1",x"72",x"32",x"c8"),
    92 => (x"6b",x"7b",x"ff",x"c3"),
    93 => (x"71",x"31",x"c8",x"4a"),
    94 => (x"7b",x"ff",x"c3",x"b2"),
    95 => (x"32",x"c8",x"49",x"6b"),
    96 => (x"48",x"71",x"b1",x"72"),
    97 => (x"4f",x"26",x"4b",x"26"),
    98 => (x"5c",x"5b",x"5e",x"0e"),
    99 => (x"4d",x"71",x"0e",x"5d"),
   100 => (x"75",x"4c",x"d4",x"ff"),
   101 => (x"98",x"ff",x"c3",x"48"),
   102 => (x"d6",x"c2",x"7c",x"70"),
   103 => (x"c8",x"05",x"bf",x"c4"),
   104 => (x"48",x"66",x"d0",x"87"),
   105 => (x"a6",x"d4",x"30",x"c9"),
   106 => (x"49",x"66",x"d0",x"58"),
   107 => (x"48",x"71",x"29",x"d8"),
   108 => (x"70",x"98",x"ff",x"c3"),
   109 => (x"49",x"66",x"d0",x"7c"),
   110 => (x"48",x"71",x"29",x"d0"),
   111 => (x"70",x"98",x"ff",x"c3"),
   112 => (x"49",x"66",x"d0",x"7c"),
   113 => (x"48",x"71",x"29",x"c8"),
   114 => (x"70",x"98",x"ff",x"c3"),
   115 => (x"48",x"66",x"d0",x"7c"),
   116 => (x"70",x"98",x"ff",x"c3"),
   117 => (x"d0",x"49",x"75",x"7c"),
   118 => (x"c3",x"48",x"71",x"29"),
   119 => (x"7c",x"70",x"98",x"ff"),
   120 => (x"f0",x"c9",x"4b",x"6c"),
   121 => (x"ff",x"c3",x"4a",x"ff"),
   122 => (x"87",x"cf",x"05",x"ab"),
   123 => (x"6c",x"7c",x"71",x"49"),
   124 => (x"02",x"8a",x"c1",x"4b"),
   125 => (x"ab",x"71",x"87",x"c5"),
   126 => (x"73",x"87",x"f2",x"02"),
   127 => (x"26",x"4d",x"26",x"48"),
   128 => (x"26",x"4b",x"26",x"4c"),
   129 => (x"49",x"c0",x"1e",x"4f"),
   130 => (x"c3",x"48",x"d4",x"ff"),
   131 => (x"81",x"c1",x"78",x"ff"),
   132 => (x"a9",x"b7",x"c8",x"c3"),
   133 => (x"26",x"87",x"f1",x"04"),
   134 => (x"5b",x"5e",x"0e",x"4f"),
   135 => (x"c0",x"0e",x"5d",x"5c"),
   136 => (x"f7",x"c1",x"f0",x"ff"),
   137 => (x"c0",x"c0",x"c1",x"4d"),
   138 => (x"4b",x"c0",x"c0",x"c0"),
   139 => (x"c4",x"87",x"d6",x"ff"),
   140 => (x"c0",x"4c",x"df",x"f8"),
   141 => (x"fd",x"49",x"75",x"1e"),
   142 => (x"86",x"c4",x"87",x"ce"),
   143 => (x"c0",x"05",x"a8",x"c1"),
   144 => (x"d4",x"ff",x"87",x"e5"),
   145 => (x"78",x"ff",x"c3",x"48"),
   146 => (x"e1",x"c0",x"1e",x"73"),
   147 => (x"49",x"e9",x"c1",x"f0"),
   148 => (x"c4",x"87",x"f5",x"fc"),
   149 => (x"05",x"98",x"70",x"86"),
   150 => (x"d4",x"ff",x"87",x"ca"),
   151 => (x"78",x"ff",x"c3",x"48"),
   152 => (x"87",x"cb",x"48",x"c1"),
   153 => (x"c1",x"87",x"de",x"fe"),
   154 => (x"c6",x"ff",x"05",x"8c"),
   155 => (x"26",x"48",x"c0",x"87"),
   156 => (x"26",x"4c",x"26",x"4d"),
   157 => (x"0e",x"4f",x"26",x"4b"),
   158 => (x"0e",x"5c",x"5b",x"5e"),
   159 => (x"c1",x"f0",x"ff",x"c0"),
   160 => (x"d4",x"ff",x"4c",x"c1"),
   161 => (x"78",x"ff",x"c3",x"48"),
   162 => (x"f8",x"49",x"fc",x"ca"),
   163 => (x"4b",x"d3",x"87",x"d9"),
   164 => (x"49",x"74",x"1e",x"c0"),
   165 => (x"c4",x"87",x"f1",x"fb"),
   166 => (x"05",x"98",x"70",x"86"),
   167 => (x"d4",x"ff",x"87",x"ca"),
   168 => (x"78",x"ff",x"c3",x"48"),
   169 => (x"87",x"cb",x"48",x"c1"),
   170 => (x"c1",x"87",x"da",x"fd"),
   171 => (x"df",x"ff",x"05",x"8b"),
   172 => (x"26",x"48",x"c0",x"87"),
   173 => (x"26",x"4b",x"26",x"4c"),
   174 => (x"00",x"00",x"00",x"4f"),
   175 => (x"00",x"44",x"4d",x"43"),
   176 => (x"43",x"48",x"44",x"53"),
   177 => (x"69",x"61",x"66",x"20"),
   178 => (x"00",x"0a",x"21",x"6c"),
   179 => (x"52",x"52",x"45",x"49"),
   180 => (x"00",x"00",x"00",x"00"),
   181 => (x"00",x"49",x"50",x"53"),
   182 => (x"74",x"69",x"72",x"57"),
   183 => (x"61",x"66",x"20",x"65"),
   184 => (x"64",x"65",x"6c",x"69"),
   185 => (x"5e",x"0e",x"00",x"0a"),
   186 => (x"0e",x"5d",x"5c",x"5b"),
   187 => (x"ff",x"4d",x"ff",x"c3"),
   188 => (x"d0",x"fc",x"4b",x"d4"),
   189 => (x"1e",x"ea",x"c6",x"87"),
   190 => (x"c1",x"f0",x"e1",x"c0"),
   191 => (x"c7",x"fa",x"49",x"c8"),
   192 => (x"c1",x"86",x"c4",x"87"),
   193 => (x"87",x"c8",x"02",x"a8"),
   194 => (x"c0",x"87",x"ec",x"fd"),
   195 => (x"87",x"e8",x"c1",x"48"),
   196 => (x"70",x"87",x"c9",x"f9"),
   197 => (x"ff",x"ff",x"cf",x"49"),
   198 => (x"a9",x"ea",x"c6",x"99"),
   199 => (x"fd",x"87",x"c8",x"02"),
   200 => (x"48",x"c0",x"87",x"d5"),
   201 => (x"75",x"87",x"d1",x"c1"),
   202 => (x"4c",x"f1",x"c0",x"7b"),
   203 => (x"70",x"87",x"ea",x"fb"),
   204 => (x"ec",x"c0",x"02",x"98"),
   205 => (x"c0",x"1e",x"c0",x"87"),
   206 => (x"fa",x"c1",x"f0",x"ff"),
   207 => (x"87",x"c8",x"f9",x"49"),
   208 => (x"98",x"70",x"86",x"c4"),
   209 => (x"75",x"87",x"da",x"05"),
   210 => (x"75",x"49",x"6b",x"7b"),
   211 => (x"75",x"7b",x"75",x"7b"),
   212 => (x"c1",x"7b",x"75",x"7b"),
   213 => (x"c4",x"02",x"99",x"c0"),
   214 => (x"db",x"48",x"c1",x"87"),
   215 => (x"d7",x"48",x"c0",x"87"),
   216 => (x"05",x"ac",x"c2",x"87"),
   217 => (x"c0",x"cb",x"87",x"ca"),
   218 => (x"87",x"fb",x"f4",x"49"),
   219 => (x"87",x"c8",x"48",x"c0"),
   220 => (x"fe",x"05",x"8c",x"c1"),
   221 => (x"48",x"c0",x"87",x"f6"),
   222 => (x"4c",x"26",x"4d",x"26"),
   223 => (x"4f",x"26",x"4b",x"26"),
   224 => (x"5c",x"5b",x"5e",x"0e"),
   225 => (x"d0",x"ff",x"0e",x"5d"),
   226 => (x"d0",x"e5",x"c0",x"4d"),
   227 => (x"c2",x"4c",x"c0",x"c1"),
   228 => (x"c1",x"48",x"c4",x"d6"),
   229 => (x"49",x"d4",x"cb",x"78"),
   230 => (x"c7",x"87",x"cc",x"f4"),
   231 => (x"f9",x"7d",x"c2",x"4b"),
   232 => (x"7d",x"c3",x"87",x"e3"),
   233 => (x"49",x"74",x"1e",x"c0"),
   234 => (x"c4",x"87",x"dd",x"f7"),
   235 => (x"05",x"a8",x"c1",x"86"),
   236 => (x"c2",x"4b",x"87",x"c1"),
   237 => (x"87",x"cb",x"05",x"ab"),
   238 => (x"f3",x"49",x"cc",x"cb"),
   239 => (x"48",x"c0",x"87",x"e9"),
   240 => (x"c1",x"87",x"f6",x"c0"),
   241 => (x"d4",x"ff",x"05",x"8b"),
   242 => (x"87",x"da",x"fc",x"87"),
   243 => (x"58",x"c8",x"d6",x"c2"),
   244 => (x"cd",x"05",x"98",x"70"),
   245 => (x"c0",x"1e",x"c1",x"87"),
   246 => (x"d0",x"c1",x"f0",x"ff"),
   247 => (x"87",x"e8",x"f6",x"49"),
   248 => (x"d4",x"ff",x"86",x"c4"),
   249 => (x"78",x"ff",x"c3",x"48"),
   250 => (x"c2",x"87",x"c3",x"c3"),
   251 => (x"c2",x"58",x"cc",x"d6"),
   252 => (x"48",x"d4",x"ff",x"7d"),
   253 => (x"c1",x"78",x"ff",x"c3"),
   254 => (x"26",x"4d",x"26",x"48"),
   255 => (x"26",x"4b",x"26",x"4c"),
   256 => (x"5b",x"5e",x"0e",x"4f"),
   257 => (x"fc",x"0e",x"5d",x"5c"),
   258 => (x"ff",x"4b",x"71",x"86"),
   259 => (x"7e",x"c0",x"4c",x"d4"),
   260 => (x"df",x"cd",x"ee",x"c5"),
   261 => (x"7c",x"ff",x"c3",x"4a"),
   262 => (x"fe",x"c3",x"48",x"6c"),
   263 => (x"f8",x"c0",x"05",x"a8"),
   264 => (x"73",x"4d",x"74",x"87"),
   265 => (x"87",x"cc",x"02",x"9b"),
   266 => (x"73",x"1e",x"66",x"d4"),
   267 => (x"87",x"c3",x"f4",x"49"),
   268 => (x"87",x"d4",x"86",x"c4"),
   269 => (x"c4",x"48",x"d0",x"ff"),
   270 => (x"66",x"d4",x"78",x"d1"),
   271 => (x"7d",x"ff",x"c3",x"4a"),
   272 => (x"f8",x"05",x"8a",x"c1"),
   273 => (x"5a",x"a6",x"d8",x"87"),
   274 => (x"7c",x"7c",x"ff",x"c3"),
   275 => (x"c5",x"05",x"9b",x"73"),
   276 => (x"48",x"d0",x"ff",x"87"),
   277 => (x"4a",x"c1",x"78",x"d0"),
   278 => (x"05",x"8a",x"c1",x"7e"),
   279 => (x"6e",x"87",x"f6",x"fe"),
   280 => (x"26",x"8e",x"fc",x"48"),
   281 => (x"26",x"4c",x"26",x"4d"),
   282 => (x"1e",x"4f",x"26",x"4b"),
   283 => (x"4a",x"71",x"1e",x"73"),
   284 => (x"d4",x"ff",x"4b",x"c0"),
   285 => (x"78",x"ff",x"c3",x"48"),
   286 => (x"c4",x"48",x"d0",x"ff"),
   287 => (x"d4",x"ff",x"78",x"c3"),
   288 => (x"78",x"ff",x"c3",x"48"),
   289 => (x"ff",x"c0",x"1e",x"72"),
   290 => (x"49",x"d1",x"c1",x"f0"),
   291 => (x"c4",x"87",x"f9",x"f3"),
   292 => (x"05",x"98",x"70",x"86"),
   293 => (x"c0",x"c8",x"87",x"d2"),
   294 => (x"49",x"66",x"cc",x"1e"),
   295 => (x"c4",x"87",x"e2",x"fd"),
   296 => (x"ff",x"4b",x"70",x"86"),
   297 => (x"78",x"c2",x"48",x"d0"),
   298 => (x"4b",x"26",x"48",x"73"),
   299 => (x"5e",x"0e",x"4f",x"26"),
   300 => (x"0e",x"5d",x"5c",x"5b"),
   301 => (x"ff",x"c0",x"1e",x"c0"),
   302 => (x"49",x"c9",x"c1",x"f0"),
   303 => (x"d2",x"87",x"c9",x"f3"),
   304 => (x"d4",x"d6",x"c2",x"1e"),
   305 => (x"87",x"f9",x"fc",x"49"),
   306 => (x"4c",x"c0",x"86",x"c8"),
   307 => (x"b7",x"d2",x"84",x"c1"),
   308 => (x"87",x"f8",x"04",x"ac"),
   309 => (x"97",x"d4",x"d6",x"c2"),
   310 => (x"c0",x"c3",x"49",x"bf"),
   311 => (x"a9",x"c0",x"c1",x"99"),
   312 => (x"87",x"e7",x"c0",x"05"),
   313 => (x"97",x"db",x"d6",x"c2"),
   314 => (x"31",x"d0",x"49",x"bf"),
   315 => (x"97",x"dc",x"d6",x"c2"),
   316 => (x"32",x"c8",x"4a",x"bf"),
   317 => (x"d6",x"c2",x"b1",x"72"),
   318 => (x"4a",x"bf",x"97",x"dd"),
   319 => (x"cf",x"4c",x"71",x"b1"),
   320 => (x"9c",x"ff",x"ff",x"ff"),
   321 => (x"34",x"ca",x"84",x"c1"),
   322 => (x"c2",x"87",x"e7",x"c1"),
   323 => (x"bf",x"97",x"dd",x"d6"),
   324 => (x"c6",x"31",x"c1",x"49"),
   325 => (x"de",x"d6",x"c2",x"99"),
   326 => (x"c7",x"4a",x"bf",x"97"),
   327 => (x"b1",x"72",x"2a",x"b7"),
   328 => (x"97",x"d9",x"d6",x"c2"),
   329 => (x"cf",x"4d",x"4a",x"bf"),
   330 => (x"da",x"d6",x"c2",x"9d"),
   331 => (x"c3",x"4a",x"bf",x"97"),
   332 => (x"c2",x"32",x"ca",x"9a"),
   333 => (x"bf",x"97",x"db",x"d6"),
   334 => (x"73",x"33",x"c2",x"4b"),
   335 => (x"dc",x"d6",x"c2",x"b2"),
   336 => (x"c3",x"4b",x"bf",x"97"),
   337 => (x"b7",x"c6",x"9b",x"c0"),
   338 => (x"c2",x"b2",x"73",x"2b"),
   339 => (x"71",x"48",x"c1",x"81"),
   340 => (x"c1",x"49",x"70",x"30"),
   341 => (x"70",x"30",x"75",x"48"),
   342 => (x"c1",x"4c",x"72",x"4d"),
   343 => (x"c8",x"94",x"71",x"84"),
   344 => (x"06",x"ad",x"b7",x"c0"),
   345 => (x"34",x"c1",x"87",x"cc"),
   346 => (x"c0",x"c8",x"2d",x"b7"),
   347 => (x"ff",x"01",x"ad",x"b7"),
   348 => (x"48",x"74",x"87",x"f4"),
   349 => (x"4c",x"26",x"4d",x"26"),
   350 => (x"4f",x"26",x"4b",x"26"),
   351 => (x"5c",x"5b",x"5e",x"0e"),
   352 => (x"86",x"f8",x"0e",x"5d"),
   353 => (x"48",x"fc",x"de",x"c2"),
   354 => (x"d6",x"c2",x"78",x"c0"),
   355 => (x"49",x"c0",x"1e",x"f4"),
   356 => (x"c4",x"87",x"d8",x"fb"),
   357 => (x"05",x"98",x"70",x"86"),
   358 => (x"48",x"c0",x"87",x"c5"),
   359 => (x"c0",x"87",x"f1",x"c8"),
   360 => (x"c2",x"7e",x"c1",x"4d"),
   361 => (x"df",x"4a",x"ea",x"d7"),
   362 => (x"4b",x"c8",x"49",x"e8"),
   363 => (x"70",x"87",x"f7",x"ec"),
   364 => (x"87",x"c2",x"05",x"98"),
   365 => (x"d8",x"c2",x"7e",x"c0"),
   366 => (x"f4",x"df",x"4a",x"c6"),
   367 => (x"ec",x"4b",x"c8",x"49"),
   368 => (x"98",x"70",x"87",x"e4"),
   369 => (x"c0",x"87",x"c2",x"05"),
   370 => (x"c0",x"02",x"6e",x"7e"),
   371 => (x"dd",x"c2",x"87",x"fd"),
   372 => (x"c2",x"4d",x"bf",x"fa"),
   373 => (x"bf",x"9f",x"f2",x"de"),
   374 => (x"d6",x"c5",x"48",x"7e"),
   375 => (x"c7",x"05",x"a8",x"ea"),
   376 => (x"fa",x"dd",x"c2",x"87"),
   377 => (x"87",x"ce",x"4d",x"bf"),
   378 => (x"e9",x"ca",x"48",x"6e"),
   379 => (x"c5",x"02",x"a8",x"d5"),
   380 => (x"c7",x"48",x"c0",x"87"),
   381 => (x"d6",x"c2",x"87",x"da"),
   382 => (x"49",x"75",x"1e",x"f4"),
   383 => (x"c4",x"87",x"ec",x"f9"),
   384 => (x"05",x"98",x"70",x"86"),
   385 => (x"48",x"c0",x"87",x"c5"),
   386 => (x"c2",x"87",x"c5",x"c7"),
   387 => (x"c0",x"4a",x"c6",x"d8"),
   388 => (x"c8",x"49",x"c0",x"e0"),
   389 => (x"87",x"ce",x"eb",x"4b"),
   390 => (x"c8",x"05",x"98",x"70"),
   391 => (x"fc",x"de",x"c2",x"87"),
   392 => (x"d7",x"78",x"c1",x"48"),
   393 => (x"ea",x"d7",x"c2",x"87"),
   394 => (x"cc",x"e0",x"c0",x"4a"),
   395 => (x"ea",x"4b",x"c8",x"49"),
   396 => (x"98",x"70",x"87",x"f4"),
   397 => (x"c0",x"87",x"c5",x"02"),
   398 => (x"87",x"d4",x"c6",x"48"),
   399 => (x"97",x"f2",x"de",x"c2"),
   400 => (x"d5",x"c1",x"49",x"bf"),
   401 => (x"87",x"cd",x"05",x"a9"),
   402 => (x"97",x"f3",x"de",x"c2"),
   403 => (x"ea",x"c2",x"49",x"bf"),
   404 => (x"c5",x"c0",x"02",x"a9"),
   405 => (x"c5",x"48",x"c0",x"87"),
   406 => (x"d6",x"c2",x"87",x"f6"),
   407 => (x"7e",x"bf",x"97",x"f4"),
   408 => (x"a8",x"e9",x"c3",x"48"),
   409 => (x"87",x"ce",x"c0",x"02"),
   410 => (x"eb",x"c3",x"48",x"6e"),
   411 => (x"c5",x"c0",x"02",x"a8"),
   412 => (x"c5",x"48",x"c0",x"87"),
   413 => (x"d6",x"c2",x"87",x"da"),
   414 => (x"49",x"bf",x"97",x"ff"),
   415 => (x"cc",x"c0",x"05",x"99"),
   416 => (x"c0",x"d7",x"c2",x"87"),
   417 => (x"c2",x"49",x"bf",x"97"),
   418 => (x"c5",x"c0",x"02",x"a9"),
   419 => (x"c4",x"48",x"c0",x"87"),
   420 => (x"d7",x"c2",x"87",x"fe"),
   421 => (x"48",x"bf",x"97",x"c1"),
   422 => (x"58",x"f8",x"de",x"c2"),
   423 => (x"c1",x"48",x"4c",x"70"),
   424 => (x"fc",x"de",x"c2",x"88"),
   425 => (x"c2",x"d7",x"c2",x"58"),
   426 => (x"75",x"49",x"bf",x"97"),
   427 => (x"c3",x"d7",x"c2",x"81"),
   428 => (x"c8",x"4a",x"bf",x"97"),
   429 => (x"7e",x"a1",x"72",x"32"),
   430 => (x"48",x"cc",x"e3",x"c2"),
   431 => (x"d7",x"c2",x"78",x"6e"),
   432 => (x"48",x"bf",x"97",x"c4"),
   433 => (x"c2",x"58",x"a6",x"c8"),
   434 => (x"02",x"bf",x"fc",x"de"),
   435 => (x"c2",x"87",x"cc",x"c2"),
   436 => (x"df",x"4a",x"c6",x"d8"),
   437 => (x"4b",x"c8",x"49",x"dc"),
   438 => (x"70",x"87",x"cb",x"e8"),
   439 => (x"c5",x"c0",x"02",x"98"),
   440 => (x"c3",x"48",x"c0",x"87"),
   441 => (x"de",x"c2",x"87",x"ea"),
   442 => (x"c2",x"4c",x"bf",x"f4"),
   443 => (x"c2",x"5c",x"e0",x"e3"),
   444 => (x"bf",x"97",x"d9",x"d7"),
   445 => (x"c2",x"31",x"c8",x"49"),
   446 => (x"bf",x"97",x"d8",x"d7"),
   447 => (x"c2",x"49",x"a1",x"4a"),
   448 => (x"bf",x"97",x"da",x"d7"),
   449 => (x"72",x"32",x"d0",x"4a"),
   450 => (x"d7",x"c2",x"49",x"a1"),
   451 => (x"4a",x"bf",x"97",x"db"),
   452 => (x"a1",x"72",x"32",x"d8"),
   453 => (x"91",x"66",x"c4",x"49"),
   454 => (x"bf",x"cc",x"e3",x"c2"),
   455 => (x"d4",x"e3",x"c2",x"81"),
   456 => (x"e1",x"d7",x"c2",x"59"),
   457 => (x"c8",x"4a",x"bf",x"97"),
   458 => (x"e0",x"d7",x"c2",x"32"),
   459 => (x"a2",x"4b",x"bf",x"97"),
   460 => (x"e2",x"d7",x"c2",x"4a"),
   461 => (x"d0",x"4b",x"bf",x"97"),
   462 => (x"4a",x"a2",x"73",x"33"),
   463 => (x"97",x"e3",x"d7",x"c2"),
   464 => (x"9b",x"cf",x"4b",x"bf"),
   465 => (x"a2",x"73",x"33",x"d8"),
   466 => (x"d8",x"e3",x"c2",x"4a"),
   467 => (x"74",x"8a",x"c2",x"5a"),
   468 => (x"d8",x"e3",x"c2",x"92"),
   469 => (x"78",x"a1",x"72",x"48"),
   470 => (x"c2",x"87",x"c1",x"c1"),
   471 => (x"bf",x"97",x"c6",x"d7"),
   472 => (x"c2",x"31",x"c8",x"49"),
   473 => (x"bf",x"97",x"c5",x"d7"),
   474 => (x"c5",x"49",x"a1",x"4a"),
   475 => (x"81",x"ff",x"c7",x"31"),
   476 => (x"e3",x"c2",x"29",x"c9"),
   477 => (x"d7",x"c2",x"59",x"e0"),
   478 => (x"4a",x"bf",x"97",x"cb"),
   479 => (x"d7",x"c2",x"32",x"c8"),
   480 => (x"4b",x"bf",x"97",x"ca"),
   481 => (x"66",x"c4",x"4a",x"a2"),
   482 => (x"c2",x"82",x"6e",x"92"),
   483 => (x"c2",x"5a",x"dc",x"e3"),
   484 => (x"c0",x"48",x"d4",x"e3"),
   485 => (x"d0",x"e3",x"c2",x"78"),
   486 => (x"78",x"a1",x"72",x"48"),
   487 => (x"48",x"e0",x"e3",x"c2"),
   488 => (x"bf",x"d4",x"e3",x"c2"),
   489 => (x"e4",x"e3",x"c2",x"78"),
   490 => (x"d8",x"e3",x"c2",x"48"),
   491 => (x"de",x"c2",x"78",x"bf"),
   492 => (x"c0",x"02",x"bf",x"fc"),
   493 => (x"48",x"74",x"87",x"c9"),
   494 => (x"7e",x"70",x"30",x"c4"),
   495 => (x"c2",x"87",x"c9",x"c0"),
   496 => (x"48",x"bf",x"dc",x"e3"),
   497 => (x"7e",x"70",x"30",x"c4"),
   498 => (x"48",x"c0",x"df",x"c2"),
   499 => (x"48",x"c1",x"78",x"6e"),
   500 => (x"4d",x"26",x"8e",x"f8"),
   501 => (x"4b",x"26",x"4c",x"26"),
   502 => (x"00",x"00",x"4f",x"26"),
   503 => (x"33",x"54",x"41",x"46"),
   504 => (x"20",x"20",x"20",x"32"),
   505 => (x"00",x"00",x"00",x"00"),
   506 => (x"31",x"54",x"41",x"46"),
   507 => (x"20",x"20",x"20",x"36"),
   508 => (x"00",x"00",x"00",x"00"),
   509 => (x"33",x"54",x"41",x"46"),
   510 => (x"20",x"20",x"20",x"32"),
   511 => (x"00",x"00",x"00",x"00"),
   512 => (x"33",x"54",x"41",x"46"),
   513 => (x"20",x"20",x"20",x"32"),
   514 => (x"00",x"00",x"00",x"00"),
   515 => (x"31",x"54",x"41",x"46"),
   516 => (x"20",x"20",x"20",x"36"),
   517 => (x"00",x"00",x"00",x"00"),
   518 => (x"20",x"20",x"2e",x"2e"),
   519 => (x"20",x"20",x"20",x"20"),
   520 => (x"00",x"20",x"20",x"20"),
   521 => (x"5c",x"5b",x"5e",x"0e"),
   522 => (x"4a",x"71",x"0e",x"5d"),
   523 => (x"bf",x"fc",x"de",x"c2"),
   524 => (x"72",x"87",x"cb",x"02"),
   525 => (x"72",x"2b",x"c7",x"4b"),
   526 => (x"9d",x"ff",x"c1",x"4d"),
   527 => (x"4b",x"72",x"87",x"c9"),
   528 => (x"4d",x"72",x"2b",x"c8"),
   529 => (x"c2",x"9d",x"ff",x"c3"),
   530 => (x"83",x"bf",x"cc",x"e3"),
   531 => (x"bf",x"c4",x"f2",x"c0"),
   532 => (x"87",x"d9",x"02",x"ab"),
   533 => (x"5b",x"c8",x"f2",x"c0"),
   534 => (x"1e",x"f4",x"d6",x"c2"),
   535 => (x"ca",x"f0",x"49",x"73"),
   536 => (x"70",x"86",x"c4",x"87"),
   537 => (x"87",x"c5",x"05",x"98"),
   538 => (x"e6",x"c0",x"48",x"c0"),
   539 => (x"fc",x"de",x"c2",x"87"),
   540 => (x"87",x"d2",x"02",x"bf"),
   541 => (x"91",x"c4",x"49",x"75"),
   542 => (x"81",x"f4",x"d6",x"c2"),
   543 => (x"ff",x"cf",x"4c",x"69"),
   544 => (x"9c",x"ff",x"ff",x"ff"),
   545 => (x"49",x"75",x"87",x"cb"),
   546 => (x"d6",x"c2",x"91",x"c2"),
   547 => (x"69",x"9f",x"81",x"f4"),
   548 => (x"26",x"48",x"74",x"4c"),
   549 => (x"26",x"4c",x"26",x"4d"),
   550 => (x"0e",x"4f",x"26",x"4b"),
   551 => (x"5d",x"5c",x"5b",x"5e"),
   552 => (x"cc",x"86",x"f4",x"0e"),
   553 => (x"66",x"c8",x"59",x"a6"),
   554 => (x"70",x"80",x"c8",x"48"),
   555 => (x"78",x"c0",x"48",x"7e"),
   556 => (x"49",x"49",x"c1",x"1e"),
   557 => (x"c4",x"87",x"d3",x"c7"),
   558 => (x"9c",x"4c",x"70",x"86"),
   559 => (x"87",x"fa",x"c0",x"02"),
   560 => (x"4a",x"c4",x"df",x"c2"),
   561 => (x"e0",x"49",x"66",x"dc"),
   562 => (x"98",x"70",x"87",x"c1"),
   563 => (x"87",x"ea",x"c0",x"02"),
   564 => (x"66",x"dc",x"4a",x"74"),
   565 => (x"e0",x"4b",x"cb",x"49"),
   566 => (x"98",x"70",x"87",x"e6"),
   567 => (x"c0",x"87",x"db",x"02"),
   568 => (x"02",x"9c",x"74",x"1e"),
   569 => (x"4d",x"c0",x"87",x"c4"),
   570 => (x"4d",x"c1",x"87",x"c2"),
   571 => (x"d9",x"c6",x"49",x"75"),
   572 => (x"70",x"86",x"c4",x"87"),
   573 => (x"ff",x"05",x"9c",x"4c"),
   574 => (x"9c",x"74",x"87",x"c6"),
   575 => (x"87",x"d7",x"c1",x"02"),
   576 => (x"6e",x"49",x"a4",x"dc"),
   577 => (x"da",x"78",x"69",x"48"),
   578 => (x"66",x"c8",x"49",x"a4"),
   579 => (x"c8",x"80",x"c4",x"48"),
   580 => (x"69",x"9f",x"58",x"a6"),
   581 => (x"08",x"66",x"c4",x"48"),
   582 => (x"fc",x"de",x"c2",x"78"),
   583 => (x"87",x"d2",x"02",x"bf"),
   584 => (x"9f",x"49",x"a4",x"d4"),
   585 => (x"ff",x"c0",x"49",x"69"),
   586 => (x"48",x"71",x"99",x"ff"),
   587 => (x"7e",x"70",x"30",x"d0"),
   588 => (x"7e",x"c0",x"87",x"c2"),
   589 => (x"66",x"c4",x"48",x"6e"),
   590 => (x"66",x"c4",x"80",x"bf"),
   591 => (x"66",x"c8",x"78",x"08"),
   592 => (x"c8",x"78",x"c0",x"48"),
   593 => (x"81",x"cc",x"49",x"66"),
   594 => (x"79",x"bf",x"66",x"c4"),
   595 => (x"d0",x"49",x"66",x"c8"),
   596 => (x"c1",x"79",x"c0",x"81"),
   597 => (x"c0",x"87",x"c2",x"48"),
   598 => (x"26",x"8e",x"f4",x"48"),
   599 => (x"26",x"4c",x"26",x"4d"),
   600 => (x"0e",x"4f",x"26",x"4b"),
   601 => (x"5d",x"5c",x"5b",x"5e"),
   602 => (x"d0",x"4c",x"71",x"0e"),
   603 => (x"6c",x"4a",x"4d",x"66"),
   604 => (x"4d",x"a1",x"72",x"49"),
   605 => (x"f8",x"de",x"c2",x"b9"),
   606 => (x"ba",x"ff",x"4a",x"bf"),
   607 => (x"99",x"71",x"99",x"72"),
   608 => (x"87",x"e4",x"c0",x"02"),
   609 => (x"6b",x"4b",x"a4",x"c4"),
   610 => (x"87",x"d8",x"fa",x"49"),
   611 => (x"de",x"c2",x"7b",x"70"),
   612 => (x"6c",x"49",x"bf",x"f4"),
   613 => (x"75",x"7c",x"71",x"81"),
   614 => (x"f8",x"de",x"c2",x"b9"),
   615 => (x"ba",x"ff",x"4a",x"bf"),
   616 => (x"99",x"71",x"99",x"72"),
   617 => (x"87",x"dc",x"ff",x"05"),
   618 => (x"4d",x"26",x"7c",x"75"),
   619 => (x"4b",x"26",x"4c",x"26"),
   620 => (x"73",x"1e",x"4f",x"26"),
   621 => (x"c2",x"4b",x"71",x"1e"),
   622 => (x"49",x"bf",x"d0",x"e3"),
   623 => (x"6a",x"4a",x"a3",x"c4"),
   624 => (x"c2",x"8a",x"c2",x"4a"),
   625 => (x"92",x"bf",x"f4",x"de"),
   626 => (x"c2",x"49",x"a1",x"72"),
   627 => (x"4a",x"bf",x"f8",x"de"),
   628 => (x"a1",x"72",x"9a",x"6b"),
   629 => (x"c8",x"f2",x"c0",x"49"),
   630 => (x"1e",x"66",x"c8",x"59"),
   631 => (x"87",x"cb",x"ea",x"71"),
   632 => (x"98",x"70",x"86",x"c4"),
   633 => (x"c0",x"87",x"c4",x"05"),
   634 => (x"c1",x"87",x"c2",x"48"),
   635 => (x"26",x"4b",x"26",x"48"),
   636 => (x"1e",x"73",x"1e",x"4f"),
   637 => (x"02",x"9b",x"4b",x"71"),
   638 => (x"c2",x"87",x"e4",x"c0"),
   639 => (x"73",x"5b",x"e4",x"e3"),
   640 => (x"c2",x"8a",x"c2",x"4a"),
   641 => (x"49",x"bf",x"f4",x"de"),
   642 => (x"d0",x"e3",x"c2",x"92"),
   643 => (x"80",x"72",x"48",x"bf"),
   644 => (x"58",x"e8",x"e3",x"c2"),
   645 => (x"30",x"c4",x"48",x"71"),
   646 => (x"58",x"c4",x"df",x"c2"),
   647 => (x"c2",x"87",x"ed",x"c0"),
   648 => (x"c2",x"48",x"e0",x"e3"),
   649 => (x"78",x"bf",x"d4",x"e3"),
   650 => (x"48",x"e4",x"e3",x"c2"),
   651 => (x"bf",x"d8",x"e3",x"c2"),
   652 => (x"fc",x"de",x"c2",x"78"),
   653 => (x"87",x"c9",x"02",x"bf"),
   654 => (x"bf",x"f4",x"de",x"c2"),
   655 => (x"c7",x"31",x"c4",x"49"),
   656 => (x"dc",x"e3",x"c2",x"87"),
   657 => (x"31",x"c4",x"49",x"bf"),
   658 => (x"59",x"c4",x"df",x"c2"),
   659 => (x"4f",x"26",x"4b",x"26"),
   660 => (x"5c",x"5b",x"5e",x"0e"),
   661 => (x"c0",x"4a",x"71",x"0e"),
   662 => (x"02",x"9a",x"72",x"4b"),
   663 => (x"da",x"87",x"e0",x"c0"),
   664 => (x"69",x"9f",x"49",x"a2"),
   665 => (x"fc",x"de",x"c2",x"4b"),
   666 => (x"87",x"cf",x"02",x"bf"),
   667 => (x"9f",x"49",x"a2",x"d4"),
   668 => (x"c0",x"4c",x"49",x"69"),
   669 => (x"d0",x"9c",x"ff",x"ff"),
   670 => (x"c0",x"87",x"c2",x"34"),
   671 => (x"73",x"b3",x"74",x"4c"),
   672 => (x"87",x"ed",x"fd",x"49"),
   673 => (x"4b",x"26",x"4c",x"26"),
   674 => (x"5e",x"0e",x"4f",x"26"),
   675 => (x"0e",x"5d",x"5c",x"5b"),
   676 => (x"a6",x"c8",x"86",x"f0"),
   677 => (x"ff",x"ff",x"cf",x"59"),
   678 => (x"c0",x"4c",x"f8",x"ff"),
   679 => (x"02",x"66",x"c4",x"7e"),
   680 => (x"d6",x"c2",x"87",x"d8"),
   681 => (x"78",x"c0",x"48",x"f0"),
   682 => (x"48",x"e8",x"d6",x"c2"),
   683 => (x"bf",x"e4",x"e3",x"c2"),
   684 => (x"ec",x"d6",x"c2",x"78"),
   685 => (x"e0",x"e3",x"c2",x"48"),
   686 => (x"df",x"c2",x"78",x"bf"),
   687 => (x"50",x"c0",x"48",x"d1"),
   688 => (x"bf",x"c0",x"df",x"c2"),
   689 => (x"f0",x"d6",x"c2",x"49"),
   690 => (x"aa",x"71",x"4a",x"bf"),
   691 => (x"87",x"cb",x"c4",x"03"),
   692 => (x"99",x"cf",x"49",x"72"),
   693 => (x"87",x"e9",x"c0",x"05"),
   694 => (x"48",x"c4",x"f2",x"c0"),
   695 => (x"bf",x"e8",x"d6",x"c2"),
   696 => (x"f4",x"d6",x"c2",x"78"),
   697 => (x"e8",x"d6",x"c2",x"1e"),
   698 => (x"d6",x"c2",x"49",x"bf"),
   699 => (x"a1",x"c1",x"48",x"e8"),
   700 => (x"f6",x"e5",x"71",x"78"),
   701 => (x"c0",x"86",x"c4",x"87"),
   702 => (x"c2",x"48",x"c0",x"f2"),
   703 => (x"cc",x"78",x"f4",x"d6"),
   704 => (x"c0",x"f2",x"c0",x"87"),
   705 => (x"e0",x"c0",x"48",x"bf"),
   706 => (x"c4",x"f2",x"c0",x"80"),
   707 => (x"f0",x"d6",x"c2",x"58"),
   708 => (x"80",x"c1",x"48",x"bf"),
   709 => (x"58",x"f4",x"d6",x"c2"),
   710 => (x"00",x"0c",x"80",x"27"),
   711 => (x"bf",x"97",x"bf",x"00"),
   712 => (x"c2",x"02",x"9d",x"4d"),
   713 => (x"e5",x"c3",x"87",x"e5"),
   714 => (x"de",x"c2",x"02",x"ad"),
   715 => (x"c0",x"f2",x"c0",x"87"),
   716 => (x"a3",x"cb",x"4b",x"bf"),
   717 => (x"cf",x"4c",x"11",x"49"),
   718 => (x"d2",x"c1",x"05",x"ac"),
   719 => (x"df",x"49",x"75",x"87"),
   720 => (x"cd",x"89",x"c1",x"99"),
   721 => (x"c4",x"df",x"c2",x"91"),
   722 => (x"4a",x"a3",x"c1",x"81"),
   723 => (x"a3",x"c3",x"51",x"12"),
   724 => (x"c5",x"51",x"12",x"4a"),
   725 => (x"51",x"12",x"4a",x"a3"),
   726 => (x"12",x"4a",x"a3",x"c7"),
   727 => (x"4a",x"a3",x"c9",x"51"),
   728 => (x"a3",x"ce",x"51",x"12"),
   729 => (x"d0",x"51",x"12",x"4a"),
   730 => (x"51",x"12",x"4a",x"a3"),
   731 => (x"12",x"4a",x"a3",x"d2"),
   732 => (x"4a",x"a3",x"d4",x"51"),
   733 => (x"a3",x"d6",x"51",x"12"),
   734 => (x"d8",x"51",x"12",x"4a"),
   735 => (x"51",x"12",x"4a",x"a3"),
   736 => (x"12",x"4a",x"a3",x"dc"),
   737 => (x"4a",x"a3",x"de",x"51"),
   738 => (x"7e",x"c1",x"51",x"12"),
   739 => (x"74",x"87",x"fc",x"c0"),
   740 => (x"05",x"99",x"c8",x"49"),
   741 => (x"74",x"87",x"ed",x"c0"),
   742 => (x"05",x"99",x"d0",x"49"),
   743 => (x"e0",x"c0",x"87",x"d3"),
   744 => (x"cc",x"c0",x"02",x"66"),
   745 => (x"c0",x"49",x"73",x"87"),
   746 => (x"70",x"0f",x"66",x"e0"),
   747 => (x"d3",x"c0",x"02",x"98"),
   748 => (x"c0",x"05",x"6e",x"87"),
   749 => (x"df",x"c2",x"87",x"c6"),
   750 => (x"50",x"c0",x"48",x"c4"),
   751 => (x"bf",x"c0",x"f2",x"c0"),
   752 => (x"87",x"e9",x"c2",x"48"),
   753 => (x"48",x"d1",x"df",x"c2"),
   754 => (x"c2",x"7e",x"50",x"c0"),
   755 => (x"49",x"bf",x"c0",x"df"),
   756 => (x"bf",x"f0",x"d6",x"c2"),
   757 => (x"04",x"aa",x"71",x"4a"),
   758 => (x"cf",x"87",x"f5",x"fb"),
   759 => (x"f8",x"ff",x"ff",x"ff"),
   760 => (x"e4",x"e3",x"c2",x"4c"),
   761 => (x"c8",x"c0",x"05",x"bf"),
   762 => (x"fc",x"de",x"c2",x"87"),
   763 => (x"fa",x"c1",x"02",x"bf"),
   764 => (x"ec",x"d6",x"c2",x"87"),
   765 => (x"eb",x"f0",x"49",x"bf"),
   766 => (x"f0",x"d6",x"c2",x"87"),
   767 => (x"48",x"a6",x"c4",x"58"),
   768 => (x"bf",x"ec",x"d6",x"c2"),
   769 => (x"fc",x"de",x"c2",x"78"),
   770 => (x"db",x"c0",x"02",x"bf"),
   771 => (x"49",x"66",x"c4",x"87"),
   772 => (x"a9",x"74",x"99",x"74"),
   773 => (x"87",x"c8",x"c0",x"02"),
   774 => (x"c0",x"48",x"a6",x"c8"),
   775 => (x"87",x"e7",x"c0",x"78"),
   776 => (x"c1",x"48",x"a6",x"c8"),
   777 => (x"87",x"df",x"c0",x"78"),
   778 => (x"cf",x"49",x"66",x"c4"),
   779 => (x"a9",x"99",x"f8",x"ff"),
   780 => (x"87",x"c8",x"c0",x"02"),
   781 => (x"c0",x"48",x"a6",x"cc"),
   782 => (x"87",x"c5",x"c0",x"78"),
   783 => (x"c1",x"48",x"a6",x"cc"),
   784 => (x"48",x"a6",x"c8",x"78"),
   785 => (x"c8",x"78",x"66",x"cc"),
   786 => (x"de",x"c0",x"05",x"66"),
   787 => (x"49",x"66",x"c4",x"87"),
   788 => (x"de",x"c2",x"89",x"c2"),
   789 => (x"c2",x"91",x"bf",x"f4"),
   790 => (x"48",x"bf",x"d0",x"e3"),
   791 => (x"d6",x"c2",x"80",x"71"),
   792 => (x"d6",x"c2",x"58",x"ec"),
   793 => (x"78",x"c0",x"48",x"f0"),
   794 => (x"c0",x"87",x"d5",x"f9"),
   795 => (x"ff",x"ff",x"cf",x"48"),
   796 => (x"f0",x"4c",x"f8",x"ff"),
   797 => (x"26",x"4d",x"26",x"8e"),
   798 => (x"26",x"4b",x"26",x"4c"),
   799 => (x"00",x"00",x"00",x"4f"),
   800 => (x"00",x"00",x"00",x"00"),
   801 => (x"ff",x"ff",x"ff",x"ff"),
   802 => (x"48",x"d4",x"ff",x"1e"),
   803 => (x"68",x"78",x"ff",x"c3"),
   804 => (x"1e",x"4f",x"26",x"48"),
   805 => (x"c3",x"48",x"d4",x"ff"),
   806 => (x"d0",x"ff",x"78",x"ff"),
   807 => (x"78",x"e1",x"c0",x"48"),
   808 => (x"d4",x"48",x"d4",x"ff"),
   809 => (x"1e",x"4f",x"26",x"78"),
   810 => (x"c0",x"48",x"d0",x"ff"),
   811 => (x"4f",x"26",x"78",x"e0"),
   812 => (x"87",x"d4",x"ff",x"1e"),
   813 => (x"02",x"99",x"49",x"70"),
   814 => (x"fb",x"c0",x"87",x"c6"),
   815 => (x"87",x"f1",x"05",x"a9"),
   816 => (x"4f",x"26",x"48",x"71"),
   817 => (x"5c",x"5b",x"5e",x"0e"),
   818 => (x"c0",x"4b",x"71",x"0e"),
   819 => (x"87",x"f8",x"fe",x"4c"),
   820 => (x"02",x"99",x"49",x"70"),
   821 => (x"c0",x"87",x"f9",x"c0"),
   822 => (x"c0",x"02",x"a9",x"ec"),
   823 => (x"fb",x"c0",x"87",x"f2"),
   824 => (x"eb",x"c0",x"02",x"a9"),
   825 => (x"b7",x"66",x"cc",x"87"),
   826 => (x"87",x"c7",x"03",x"ac"),
   827 => (x"c2",x"02",x"66",x"d0"),
   828 => (x"71",x"53",x"71",x"87"),
   829 => (x"87",x"c2",x"02",x"99"),
   830 => (x"cb",x"fe",x"84",x"c1"),
   831 => (x"99",x"49",x"70",x"87"),
   832 => (x"c0",x"87",x"cd",x"02"),
   833 => (x"c7",x"02",x"a9",x"ec"),
   834 => (x"a9",x"fb",x"c0",x"87"),
   835 => (x"87",x"d5",x"ff",x"05"),
   836 => (x"c3",x"02",x"66",x"d0"),
   837 => (x"7b",x"97",x"c0",x"87"),
   838 => (x"05",x"a9",x"ec",x"c0"),
   839 => (x"4a",x"74",x"87",x"c4"),
   840 => (x"4a",x"74",x"87",x"c5"),
   841 => (x"72",x"8a",x"0a",x"c0"),
   842 => (x"26",x"4c",x"26",x"48"),
   843 => (x"1e",x"4f",x"26",x"4b"),
   844 => (x"70",x"87",x"d5",x"fd"),
   845 => (x"f0",x"c0",x"4a",x"49"),
   846 => (x"87",x"c9",x"04",x"aa"),
   847 => (x"01",x"aa",x"f9",x"c0"),
   848 => (x"f0",x"c0",x"87",x"c3"),
   849 => (x"aa",x"c1",x"c1",x"8a"),
   850 => (x"c1",x"87",x"c9",x"04"),
   851 => (x"c3",x"01",x"aa",x"da"),
   852 => (x"8a",x"f7",x"c0",x"87"),
   853 => (x"4f",x"26",x"48",x"72"),
   854 => (x"5c",x"5b",x"5e",x"0e"),
   855 => (x"86",x"f8",x"0e",x"5d"),
   856 => (x"7e",x"c0",x"4c",x"71"),
   857 => (x"c0",x"87",x"ec",x"fc"),
   858 => (x"f8",x"f7",x"c0",x"4b"),
   859 => (x"c0",x"49",x"bf",x"97"),
   860 => (x"87",x"cf",x"04",x"a9"),
   861 => (x"c1",x"87",x"f9",x"fc"),
   862 => (x"f8",x"f7",x"c0",x"83"),
   863 => (x"ab",x"49",x"bf",x"97"),
   864 => (x"c0",x"87",x"f1",x"06"),
   865 => (x"bf",x"97",x"f8",x"f7"),
   866 => (x"fb",x"87",x"cf",x"02"),
   867 => (x"49",x"70",x"87",x"fa"),
   868 => (x"87",x"c6",x"02",x"99"),
   869 => (x"05",x"a9",x"ec",x"c0"),
   870 => (x"4b",x"c0",x"87",x"f1"),
   871 => (x"70",x"87",x"e9",x"fb"),
   872 => (x"87",x"e4",x"fb",x"4d"),
   873 => (x"fb",x"58",x"a6",x"c8"),
   874 => (x"4a",x"70",x"87",x"de"),
   875 => (x"a4",x"c8",x"83",x"c1"),
   876 => (x"49",x"69",x"97",x"49"),
   877 => (x"87",x"da",x"05",x"ad"),
   878 => (x"97",x"49",x"a4",x"c9"),
   879 => (x"66",x"c4",x"49",x"69"),
   880 => (x"87",x"ce",x"05",x"a9"),
   881 => (x"97",x"49",x"a4",x"ca"),
   882 => (x"05",x"aa",x"49",x"69"),
   883 => (x"7e",x"c1",x"87",x"c4"),
   884 => (x"ec",x"c0",x"87",x"d0"),
   885 => (x"87",x"c6",x"02",x"ad"),
   886 => (x"05",x"ad",x"fb",x"c0"),
   887 => (x"4b",x"c0",x"87",x"c4"),
   888 => (x"02",x"6e",x"7e",x"c1"),
   889 => (x"fa",x"87",x"f5",x"fe"),
   890 => (x"48",x"73",x"87",x"fd"),
   891 => (x"4d",x"26",x"8e",x"f8"),
   892 => (x"4b",x"26",x"4c",x"26"),
   893 => (x"00",x"00",x"4f",x"26"),
   894 => (x"1e",x"73",x"1e",x"00"),
   895 => (x"c8",x"4b",x"d4",x"ff"),
   896 => (x"d0",x"ff",x"4a",x"66"),
   897 => (x"78",x"c5",x"c8",x"48"),
   898 => (x"c1",x"48",x"d4",x"ff"),
   899 => (x"7b",x"11",x"78",x"d4"),
   900 => (x"f9",x"05",x"8a",x"c1"),
   901 => (x"48",x"d0",x"ff",x"87"),
   902 => (x"4b",x"26",x"78",x"c4"),
   903 => (x"5e",x"0e",x"4f",x"26"),
   904 => (x"0e",x"5d",x"5c",x"5b"),
   905 => (x"7e",x"71",x"86",x"f8"),
   906 => (x"e3",x"c2",x"1e",x"6e"),
   907 => (x"ea",x"e9",x"49",x"f4"),
   908 => (x"70",x"86",x"c4",x"87"),
   909 => (x"e4",x"c4",x"02",x"98"),
   910 => (x"cc",x"e6",x"c1",x"87"),
   911 => (x"49",x"6e",x"4c",x"bf"),
   912 => (x"c8",x"87",x"d5",x"fc"),
   913 => (x"98",x"70",x"58",x"a6"),
   914 => (x"c4",x"87",x"c5",x"05"),
   915 => (x"78",x"c1",x"48",x"a6"),
   916 => (x"c5",x"48",x"d0",x"ff"),
   917 => (x"48",x"d4",x"ff",x"78"),
   918 => (x"c4",x"78",x"d5",x"c1"),
   919 => (x"89",x"c1",x"49",x"66"),
   920 => (x"e6",x"c1",x"31",x"c6"),
   921 => (x"4a",x"bf",x"97",x"c4"),
   922 => (x"ff",x"b0",x"71",x"48"),
   923 => (x"ff",x"78",x"08",x"d4"),
   924 => (x"78",x"c4",x"48",x"d0"),
   925 => (x"97",x"f0",x"e3",x"c2"),
   926 => (x"99",x"d0",x"49",x"bf"),
   927 => (x"c5",x"87",x"dd",x"02"),
   928 => (x"48",x"d4",x"ff",x"78"),
   929 => (x"c0",x"78",x"d6",x"c1"),
   930 => (x"48",x"d4",x"ff",x"4a"),
   931 => (x"c1",x"78",x"ff",x"c3"),
   932 => (x"aa",x"e0",x"c0",x"82"),
   933 => (x"ff",x"87",x"f2",x"04"),
   934 => (x"78",x"c4",x"48",x"d0"),
   935 => (x"c3",x"48",x"d4",x"ff"),
   936 => (x"d0",x"ff",x"78",x"ff"),
   937 => (x"ff",x"78",x"c5",x"48"),
   938 => (x"d3",x"c1",x"48",x"d4"),
   939 => (x"ff",x"78",x"c1",x"78"),
   940 => (x"78",x"c4",x"48",x"d0"),
   941 => (x"06",x"ac",x"b7",x"c0"),
   942 => (x"c2",x"87",x"cb",x"c2"),
   943 => (x"4b",x"bf",x"fc",x"e3"),
   944 => (x"73",x"7e",x"74",x"8c"),
   945 => (x"dd",x"c1",x"02",x"9b"),
   946 => (x"4d",x"c0",x"c8",x"87"),
   947 => (x"ab",x"b7",x"c0",x"8b"),
   948 => (x"c8",x"87",x"c6",x"03"),
   949 => (x"c0",x"4d",x"a3",x"c0"),
   950 => (x"f0",x"e3",x"c2",x"4b"),
   951 => (x"d0",x"49",x"bf",x"97"),
   952 => (x"87",x"cf",x"02",x"99"),
   953 => (x"e3",x"c2",x"1e",x"c0"),
   954 => (x"c5",x"eb",x"49",x"f4"),
   955 => (x"70",x"86",x"c4",x"87"),
   956 => (x"c2",x"87",x"d8",x"4c"),
   957 => (x"c2",x"1e",x"f4",x"d6"),
   958 => (x"ea",x"49",x"f4",x"e3"),
   959 => (x"4c",x"70",x"87",x"f4"),
   960 => (x"d6",x"c2",x"1e",x"75"),
   961 => (x"f0",x"fb",x"49",x"f4"),
   962 => (x"74",x"86",x"c8",x"87"),
   963 => (x"87",x"c5",x"05",x"9c"),
   964 => (x"ca",x"c1",x"48",x"c0"),
   965 => (x"c2",x"1e",x"c1",x"87"),
   966 => (x"e9",x"49",x"f4",x"e3"),
   967 => (x"86",x"c4",x"87",x"c5"),
   968 => (x"fe",x"05",x"9b",x"73"),
   969 => (x"4c",x"6e",x"87",x"e3"),
   970 => (x"06",x"ac",x"b7",x"c0"),
   971 => (x"e3",x"c2",x"87",x"d1"),
   972 => (x"78",x"c0",x"48",x"f4"),
   973 => (x"78",x"c0",x"80",x"d0"),
   974 => (x"e4",x"c2",x"80",x"f4"),
   975 => (x"c0",x"78",x"bf",x"c0"),
   976 => (x"fd",x"01",x"ac",x"b7"),
   977 => (x"d0",x"ff",x"87",x"f5"),
   978 => (x"ff",x"78",x"c5",x"48"),
   979 => (x"d3",x"c1",x"48",x"d4"),
   980 => (x"ff",x"78",x"c0",x"78"),
   981 => (x"78",x"c4",x"48",x"d0"),
   982 => (x"c2",x"c0",x"48",x"c1"),
   983 => (x"f8",x"48",x"c0",x"87"),
   984 => (x"26",x"4d",x"26",x"8e"),
   985 => (x"26",x"4b",x"26",x"4c"),
   986 => (x"5b",x"5e",x"0e",x"4f"),
   987 => (x"fc",x"0e",x"5d",x"5c"),
   988 => (x"c0",x"4d",x"71",x"86"),
   989 => (x"04",x"ad",x"4c",x"4b"),
   990 => (x"c0",x"87",x"e8",x"c0"),
   991 => (x"74",x"1e",x"d8",x"f5"),
   992 => (x"87",x"c4",x"02",x"9c"),
   993 => (x"87",x"c2",x"4a",x"c0"),
   994 => (x"49",x"72",x"4a",x"c1"),
   995 => (x"c4",x"87",x"fb",x"eb"),
   996 => (x"c1",x"7e",x"70",x"86"),
   997 => (x"c2",x"05",x"6e",x"83"),
   998 => (x"c1",x"4b",x"75",x"87"),
   999 => (x"06",x"ab",x"75",x"84"),
  1000 => (x"6e",x"87",x"d8",x"ff"),
  1001 => (x"26",x"8e",x"fc",x"48"),
  1002 => (x"26",x"4c",x"26",x"4d"),
  1003 => (x"1e",x"4f",x"26",x"4b"),
  1004 => (x"66",x"c4",x"4a",x"71"),
  1005 => (x"72",x"87",x"c5",x"05"),
  1006 => (x"87",x"e2",x"f9",x"49"),
  1007 => (x"5e",x"0e",x"4f",x"26"),
  1008 => (x"0e",x"5d",x"5c",x"5b"),
  1009 => (x"4c",x"71",x"86",x"fc"),
  1010 => (x"c2",x"91",x"de",x"49"),
  1011 => (x"71",x"4d",x"e0",x"e4"),
  1012 => (x"02",x"6d",x"97",x"85"),
  1013 => (x"c2",x"87",x"dc",x"c1"),
  1014 => (x"49",x"bf",x"d0",x"e4"),
  1015 => (x"fe",x"71",x"81",x"74"),
  1016 => (x"7e",x"70",x"87",x"c7"),
  1017 => (x"c0",x"02",x"98",x"48"),
  1018 => (x"e4",x"c2",x"87",x"f2"),
  1019 => (x"4a",x"70",x"4b",x"d4"),
  1020 => (x"c4",x"ff",x"49",x"cb"),
  1021 => (x"4b",x"74",x"87",x"ed"),
  1022 => (x"e6",x"c1",x"93",x"cc"),
  1023 => (x"83",x"c4",x"83",x"d0"),
  1024 => (x"7b",x"c0",x"c1",x"c1"),
  1025 => (x"c4",x"c1",x"49",x"74"),
  1026 => (x"7b",x"75",x"87",x"ce"),
  1027 => (x"97",x"c8",x"e6",x"c1"),
  1028 => (x"c2",x"1e",x"49",x"bf"),
  1029 => (x"fe",x"49",x"d4",x"e4"),
  1030 => (x"86",x"c4",x"87",x"d5"),
  1031 => (x"c3",x"c1",x"49",x"74"),
  1032 => (x"49",x"c0",x"87",x"f6"),
  1033 => (x"87",x"d1",x"c5",x"c1"),
  1034 => (x"48",x"ec",x"e3",x"c2"),
  1035 => (x"c0",x"49",x"50",x"c0"),
  1036 => (x"fc",x"87",x"e6",x"e2"),
  1037 => (x"26",x"4d",x"26",x"8e"),
  1038 => (x"26",x"4b",x"26",x"4c"),
  1039 => (x"00",x"00",x"00",x"4f"),
  1040 => (x"64",x"61",x"6f",x"4c"),
  1041 => (x"2e",x"67",x"6e",x"69"),
  1042 => (x"00",x"00",x"2e",x"2e"),
  1043 => (x"61",x"42",x"20",x"80"),
  1044 => (x"00",x"00",x"6b",x"63"),
  1045 => (x"64",x"61",x"6f",x"4c"),
  1046 => (x"20",x"2e",x"2a",x"20"),
  1047 => (x"00",x"00",x"00",x"00"),
  1048 => (x"00",x"00",x"20",x"3a"),
  1049 => (x"61",x"42",x"20",x"80"),
  1050 => (x"00",x"00",x"6b",x"63"),
  1051 => (x"78",x"45",x"20",x"80"),
  1052 => (x"00",x"00",x"74",x"69"),
  1053 => (x"49",x"20",x"44",x"53"),
  1054 => (x"2e",x"74",x"69",x"6e"),
  1055 => (x"00",x"00",x"00",x"2e"),
  1056 => (x"00",x"00",x"4b",x"4f"),
  1057 => (x"54",x"4f",x"4f",x"42"),
  1058 => (x"20",x"20",x"20",x"20"),
  1059 => (x"00",x"4d",x"4f",x"52"),
  1060 => (x"71",x"1e",x"73",x"1e"),
  1061 => (x"e4",x"c2",x"49",x"4b"),
  1062 => (x"71",x"81",x"bf",x"d0"),
  1063 => (x"70",x"87",x"ca",x"fb"),
  1064 => (x"c4",x"02",x"9a",x"4a"),
  1065 => (x"e7",x"e6",x"49",x"87"),
  1066 => (x"d0",x"e4",x"c2",x"87"),
  1067 => (x"73",x"78",x"c0",x"48"),
  1068 => (x"87",x"fa",x"c1",x"49"),
  1069 => (x"4f",x"26",x"4b",x"26"),
  1070 => (x"71",x"1e",x"73",x"1e"),
  1071 => (x"4a",x"a3",x"c4",x"4b"),
  1072 => (x"87",x"d0",x"c1",x"02"),
  1073 => (x"dc",x"02",x"8a",x"c1"),
  1074 => (x"c0",x"02",x"8a",x"87"),
  1075 => (x"05",x"8a",x"87",x"f2"),
  1076 => (x"c2",x"87",x"d3",x"c1"),
  1077 => (x"02",x"bf",x"d0",x"e4"),
  1078 => (x"48",x"87",x"cb",x"c1"),
  1079 => (x"e4",x"c2",x"88",x"c1"),
  1080 => (x"c1",x"c1",x"58",x"d4"),
  1081 => (x"d0",x"e4",x"c2",x"87"),
  1082 => (x"89",x"c6",x"49",x"bf"),
  1083 => (x"59",x"d4",x"e4",x"c2"),
  1084 => (x"03",x"a9",x"b7",x"c0"),
  1085 => (x"c2",x"87",x"ef",x"c0"),
  1086 => (x"c0",x"48",x"d0",x"e4"),
  1087 => (x"87",x"e6",x"c0",x"78"),
  1088 => (x"bf",x"cc",x"e4",x"c2"),
  1089 => (x"c2",x"87",x"df",x"02"),
  1090 => (x"48",x"bf",x"d0",x"e4"),
  1091 => (x"e4",x"c2",x"80",x"c1"),
  1092 => (x"87",x"d2",x"58",x"d4"),
  1093 => (x"bf",x"cc",x"e4",x"c2"),
  1094 => (x"c2",x"87",x"cb",x"02"),
  1095 => (x"48",x"bf",x"d0",x"e4"),
  1096 => (x"e4",x"c2",x"80",x"c6"),
  1097 => (x"49",x"73",x"58",x"d4"),
  1098 => (x"4b",x"26",x"87",x"c4"),
  1099 => (x"5e",x"0e",x"4f",x"26"),
  1100 => (x"0e",x"5d",x"5c",x"5b"),
  1101 => (x"a6",x"d0",x"86",x"f0"),
  1102 => (x"f4",x"d6",x"c2",x"59"),
  1103 => (x"c2",x"4c",x"c0",x"4d"),
  1104 => (x"c1",x"48",x"cc",x"e4"),
  1105 => (x"48",x"a6",x"c8",x"78"),
  1106 => (x"7e",x"75",x"78",x"c0"),
  1107 => (x"bf",x"d0",x"e4",x"c2"),
  1108 => (x"06",x"a8",x"c0",x"48"),
  1109 => (x"c8",x"87",x"c0",x"c1"),
  1110 => (x"7e",x"75",x"5c",x"a6"),
  1111 => (x"48",x"f4",x"d6",x"c2"),
  1112 => (x"f2",x"c0",x"02",x"98"),
  1113 => (x"4d",x"66",x"c4",x"87"),
  1114 => (x"1e",x"d8",x"f5",x"c0"),
  1115 => (x"c4",x"02",x"66",x"cc"),
  1116 => (x"c2",x"4c",x"c0",x"87"),
  1117 => (x"74",x"4c",x"c1",x"87"),
  1118 => (x"87",x"ce",x"e4",x"49"),
  1119 => (x"7e",x"70",x"86",x"c4"),
  1120 => (x"66",x"c8",x"85",x"c1"),
  1121 => (x"cc",x"80",x"c1",x"48"),
  1122 => (x"e4",x"c2",x"58",x"a6"),
  1123 => (x"03",x"ad",x"bf",x"d0"),
  1124 => (x"05",x"6e",x"87",x"c5"),
  1125 => (x"6e",x"87",x"d1",x"ff"),
  1126 => (x"75",x"4c",x"c0",x"4d"),
  1127 => (x"dc",x"c3",x"02",x"9d"),
  1128 => (x"d8",x"f5",x"c0",x"87"),
  1129 => (x"02",x"66",x"cc",x"1e"),
  1130 => (x"a6",x"c8",x"87",x"c7"),
  1131 => (x"c5",x"78",x"c0",x"48"),
  1132 => (x"48",x"a6",x"c8",x"87"),
  1133 => (x"66",x"c8",x"78",x"c1"),
  1134 => (x"87",x"ce",x"e3",x"49"),
  1135 => (x"7e",x"70",x"86",x"c4"),
  1136 => (x"c2",x"02",x"98",x"48"),
  1137 => (x"cb",x"49",x"87",x"e4"),
  1138 => (x"49",x"69",x"97",x"81"),
  1139 => (x"c1",x"02",x"99",x"d0"),
  1140 => (x"49",x"74",x"87",x"d4"),
  1141 => (x"e6",x"c1",x"91",x"cc"),
  1142 => (x"c2",x"c1",x"81",x"d0"),
  1143 => (x"81",x"c8",x"79",x"d0"),
  1144 => (x"74",x"51",x"ff",x"c3"),
  1145 => (x"c2",x"91",x"de",x"49"),
  1146 => (x"71",x"4d",x"e0",x"e4"),
  1147 => (x"97",x"c1",x"c2",x"85"),
  1148 => (x"49",x"a5",x"c1",x"7d"),
  1149 => (x"c2",x"51",x"e0",x"c0"),
  1150 => (x"bf",x"97",x"c4",x"df"),
  1151 => (x"c1",x"87",x"d2",x"02"),
  1152 => (x"4b",x"a5",x"c2",x"84"),
  1153 => (x"4a",x"c4",x"df",x"c2"),
  1154 => (x"fc",x"fe",x"49",x"db"),
  1155 => (x"d9",x"c1",x"87",x"d5"),
  1156 => (x"49",x"a5",x"cd",x"87"),
  1157 => (x"84",x"c1",x"51",x"c0"),
  1158 => (x"6e",x"4b",x"a5",x"c2"),
  1159 => (x"fe",x"49",x"cb",x"4a"),
  1160 => (x"c1",x"87",x"c0",x"fc"),
  1161 => (x"49",x"74",x"87",x"c4"),
  1162 => (x"e6",x"c1",x"91",x"cc"),
  1163 => (x"fe",x"c0",x"81",x"d0"),
  1164 => (x"df",x"c2",x"79",x"fe"),
  1165 => (x"02",x"bf",x"97",x"c4"),
  1166 => (x"49",x"74",x"87",x"d8"),
  1167 => (x"84",x"c1",x"91",x"de"),
  1168 => (x"4b",x"e0",x"e4",x"c2"),
  1169 => (x"df",x"c2",x"83",x"71"),
  1170 => (x"49",x"dd",x"4a",x"c4"),
  1171 => (x"87",x"d3",x"fb",x"fe"),
  1172 => (x"4b",x"74",x"87",x"d8"),
  1173 => (x"e4",x"c2",x"93",x"de"),
  1174 => (x"a3",x"cb",x"83",x"e0"),
  1175 => (x"c1",x"51",x"c0",x"49"),
  1176 => (x"4a",x"6e",x"73",x"84"),
  1177 => (x"fa",x"fe",x"49",x"cb"),
  1178 => (x"66",x"c8",x"87",x"f9"),
  1179 => (x"cc",x"80",x"c1",x"48"),
  1180 => (x"ac",x"c7",x"58",x"a6"),
  1181 => (x"87",x"c5",x"c0",x"03"),
  1182 => (x"e4",x"fc",x"05",x"6e"),
  1183 => (x"03",x"ac",x"c7",x"87"),
  1184 => (x"c2",x"87",x"e4",x"c0"),
  1185 => (x"c0",x"48",x"cc",x"e4"),
  1186 => (x"cc",x"49",x"74",x"78"),
  1187 => (x"d0",x"e6",x"c1",x"91"),
  1188 => (x"fe",x"fe",x"c0",x"81"),
  1189 => (x"de",x"49",x"74",x"79"),
  1190 => (x"e0",x"e4",x"c2",x"91"),
  1191 => (x"c1",x"51",x"c0",x"81"),
  1192 => (x"04",x"ac",x"c7",x"84"),
  1193 => (x"c1",x"87",x"dc",x"ff"),
  1194 => (x"c0",x"48",x"ec",x"e7"),
  1195 => (x"c1",x"80",x"f7",x"50"),
  1196 => (x"c1",x"40",x"d4",x"cc"),
  1197 => (x"c8",x"78",x"cc",x"c1"),
  1198 => (x"f8",x"c2",x"c1",x"80"),
  1199 => (x"49",x"66",x"cc",x"78"),
  1200 => (x"87",x"d4",x"f9",x"c0"),
  1201 => (x"4d",x"26",x"8e",x"f0"),
  1202 => (x"4b",x"26",x"4c",x"26"),
  1203 => (x"73",x"1e",x"4f",x"26"),
  1204 => (x"49",x"4b",x"71",x"1e"),
  1205 => (x"e6",x"c1",x"91",x"cc"),
  1206 => (x"a1",x"c8",x"81",x"d0"),
  1207 => (x"c4",x"e6",x"c1",x"4a"),
  1208 => (x"c9",x"50",x"12",x"48"),
  1209 => (x"f7",x"c0",x"4a",x"a1"),
  1210 => (x"50",x"12",x"48",x"f8"),
  1211 => (x"e6",x"c1",x"81",x"ca"),
  1212 => (x"50",x"11",x"48",x"c8"),
  1213 => (x"97",x"c8",x"e6",x"c1"),
  1214 => (x"c0",x"1e",x"49",x"bf"),
  1215 => (x"87",x"ef",x"f2",x"49"),
  1216 => (x"e9",x"f8",x"49",x"73"),
  1217 => (x"26",x"8e",x"fc",x"87"),
  1218 => (x"1e",x"4f",x"26",x"4b"),
  1219 => (x"f9",x"c0",x"49",x"c0"),
  1220 => (x"4f",x"26",x"87",x"e7"),
  1221 => (x"49",x"4a",x"71",x"1e"),
  1222 => (x"e6",x"c1",x"91",x"cc"),
  1223 => (x"81",x"c8",x"81",x"d0"),
  1224 => (x"48",x"ec",x"e3",x"c2"),
  1225 => (x"f0",x"c0",x"50",x"11"),
  1226 => (x"f5",x"fe",x"49",x"a2"),
  1227 => (x"49",x"c0",x"87",x"de"),
  1228 => (x"26",x"87",x"e6",x"d6"),
  1229 => (x"d4",x"ff",x"1e",x"4f"),
  1230 => (x"7a",x"ff",x"c3",x"4a"),
  1231 => (x"c0",x"48",x"d0",x"ff"),
  1232 => (x"7a",x"de",x"78",x"e1"),
  1233 => (x"c8",x"48",x"7a",x"71"),
  1234 => (x"7a",x"70",x"28",x"b7"),
  1235 => (x"b7",x"d0",x"48",x"71"),
  1236 => (x"71",x"7a",x"70",x"28"),
  1237 => (x"28",x"b7",x"d8",x"48"),
  1238 => (x"d0",x"ff",x"7a",x"70"),
  1239 => (x"78",x"e0",x"c0",x"48"),
  1240 => (x"5e",x"0e",x"4f",x"26"),
  1241 => (x"0e",x"5d",x"5c",x"5b"),
  1242 => (x"4d",x"71",x"86",x"f4"),
  1243 => (x"c1",x"91",x"cc",x"49"),
  1244 => (x"c8",x"81",x"d0",x"e6"),
  1245 => (x"a1",x"ca",x"4a",x"a1"),
  1246 => (x"48",x"a6",x"c4",x"7e"),
  1247 => (x"bf",x"e8",x"e3",x"c2"),
  1248 => (x"bf",x"97",x"6e",x"78"),
  1249 => (x"4c",x"66",x"c4",x"4b"),
  1250 => (x"48",x"12",x"2c",x"73"),
  1251 => (x"70",x"58",x"a6",x"cc"),
  1252 => (x"c9",x"84",x"c1",x"9c"),
  1253 => (x"49",x"69",x"97",x"81"),
  1254 => (x"c2",x"04",x"ac",x"b7"),
  1255 => (x"6e",x"4c",x"c0",x"87"),
  1256 => (x"c8",x"4a",x"bf",x"97"),
  1257 => (x"31",x"72",x"49",x"66"),
  1258 => (x"66",x"c4",x"b9",x"ff"),
  1259 => (x"72",x"48",x"74",x"99"),
  1260 => (x"b1",x"4a",x"70",x"30"),
  1261 => (x"59",x"ec",x"e3",x"c2"),
  1262 => (x"87",x"f9",x"fd",x"71"),
  1263 => (x"e4",x"c2",x"1e",x"c7"),
  1264 => (x"c1",x"1e",x"bf",x"c8"),
  1265 => (x"c2",x"1e",x"d0",x"e6"),
  1266 => (x"bf",x"97",x"ec",x"e3"),
  1267 => (x"87",x"f4",x"c1",x"49"),
  1268 => (x"f5",x"c0",x"49",x"75"),
  1269 => (x"8e",x"e8",x"87",x"c2"),
  1270 => (x"4c",x"26",x"4d",x"26"),
  1271 => (x"4f",x"26",x"4b",x"26"),
  1272 => (x"71",x"1e",x"73",x"1e"),
  1273 => (x"f9",x"fd",x"49",x"4b"),
  1274 => (x"fd",x"49",x"73",x"87"),
  1275 => (x"4b",x"26",x"87",x"f4"),
  1276 => (x"73",x"1e",x"4f",x"26"),
  1277 => (x"c2",x"4b",x"71",x"1e"),
  1278 => (x"d6",x"02",x"4a",x"a3"),
  1279 => (x"05",x"8a",x"c1",x"87"),
  1280 => (x"c2",x"87",x"e2",x"c0"),
  1281 => (x"02",x"bf",x"c8",x"e4"),
  1282 => (x"c1",x"48",x"87",x"db"),
  1283 => (x"cc",x"e4",x"c2",x"88"),
  1284 => (x"c2",x"87",x"d2",x"58"),
  1285 => (x"02",x"bf",x"cc",x"e4"),
  1286 => (x"e4",x"c2",x"87",x"cb"),
  1287 => (x"c1",x"48",x"bf",x"c8"),
  1288 => (x"cc",x"e4",x"c2",x"80"),
  1289 => (x"c2",x"1e",x"c7",x"58"),
  1290 => (x"1e",x"bf",x"c8",x"e4"),
  1291 => (x"1e",x"d0",x"e6",x"c1"),
  1292 => (x"97",x"ec",x"e3",x"c2"),
  1293 => (x"87",x"cc",x"49",x"bf"),
  1294 => (x"f3",x"c0",x"49",x"73"),
  1295 => (x"8e",x"f4",x"87",x"da"),
  1296 => (x"4f",x"26",x"4b",x"26"),
  1297 => (x"5c",x"5b",x"5e",x"0e"),
  1298 => (x"cc",x"ff",x"0e",x"5d"),
  1299 => (x"a6",x"e4",x"c0",x"86"),
  1300 => (x"48",x"a6",x"cc",x"59"),
  1301 => (x"80",x"c4",x"78",x"c0"),
  1302 => (x"80",x"c4",x"78",x"c0"),
  1303 => (x"78",x"66",x"c8",x"c1"),
  1304 => (x"78",x"c1",x"80",x"c4"),
  1305 => (x"78",x"c1",x"80",x"c4"),
  1306 => (x"48",x"cc",x"e4",x"c2"),
  1307 => (x"e2",x"e0",x"78",x"c1"),
  1308 => (x"87",x"fc",x"e0",x"87"),
  1309 => (x"70",x"87",x"d1",x"e0"),
  1310 => (x"ac",x"fb",x"c0",x"4c"),
  1311 => (x"87",x"f3",x"c1",x"02"),
  1312 => (x"05",x"66",x"e0",x"c0"),
  1313 => (x"c1",x"87",x"e8",x"c1"),
  1314 => (x"c4",x"4a",x"66",x"c4"),
  1315 => (x"c1",x"7e",x"6a",x"82"),
  1316 => (x"6e",x"48",x"d4",x"c1"),
  1317 => (x"20",x"41",x"20",x"49"),
  1318 => (x"c1",x"51",x"10",x"41"),
  1319 => (x"c1",x"48",x"66",x"c4"),
  1320 => (x"6a",x"78",x"ce",x"cb"),
  1321 => (x"74",x"81",x"c7",x"49"),
  1322 => (x"66",x"c4",x"c1",x"51"),
  1323 => (x"c1",x"81",x"c8",x"49"),
  1324 => (x"48",x"a6",x"d8",x"51"),
  1325 => (x"c4",x"c1",x"78",x"c2"),
  1326 => (x"81",x"c9",x"49",x"66"),
  1327 => (x"c4",x"c1",x"51",x"c0"),
  1328 => (x"81",x"ca",x"49",x"66"),
  1329 => (x"1e",x"c1",x"51",x"c0"),
  1330 => (x"49",x"6a",x"1e",x"d8"),
  1331 => (x"df",x"ff",x"81",x"c8"),
  1332 => (x"86",x"c8",x"87",x"f2"),
  1333 => (x"48",x"66",x"c8",x"c1"),
  1334 => (x"c7",x"01",x"a8",x"c0"),
  1335 => (x"48",x"a6",x"d0",x"87"),
  1336 => (x"87",x"cf",x"78",x"c1"),
  1337 => (x"48",x"66",x"c8",x"c1"),
  1338 => (x"a6",x"d8",x"88",x"c1"),
  1339 => (x"ff",x"87",x"c4",x"58"),
  1340 => (x"74",x"87",x"fd",x"de"),
  1341 => (x"da",x"cd",x"02",x"9c"),
  1342 => (x"48",x"66",x"d0",x"87"),
  1343 => (x"a8",x"66",x"cc",x"c1"),
  1344 => (x"87",x"cf",x"cd",x"03"),
  1345 => (x"c0",x"48",x"a6",x"c8"),
  1346 => (x"dd",x"ff",x"7e",x"78"),
  1347 => (x"4c",x"70",x"87",x"fa"),
  1348 => (x"05",x"ac",x"d0",x"c1"),
  1349 => (x"c4",x"87",x"e7",x"c2"),
  1350 => (x"78",x"6e",x"48",x"a6"),
  1351 => (x"70",x"87",x"d0",x"e0"),
  1352 => (x"66",x"cc",x"48",x"7e"),
  1353 => (x"87",x"c5",x"06",x"a8"),
  1354 => (x"6e",x"48",x"a6",x"cc"),
  1355 => (x"d7",x"dd",x"ff",x"78"),
  1356 => (x"c0",x"4c",x"70",x"87"),
  1357 => (x"c1",x"05",x"ac",x"ec"),
  1358 => (x"66",x"d0",x"87",x"ee"),
  1359 => (x"c1",x"91",x"cc",x"49"),
  1360 => (x"c4",x"81",x"66",x"c4"),
  1361 => (x"4d",x"6a",x"4a",x"a1"),
  1362 => (x"6e",x"4a",x"a1",x"c8"),
  1363 => (x"d4",x"cc",x"c1",x"52"),
  1364 => (x"f3",x"dc",x"ff",x"79"),
  1365 => (x"9c",x"4c",x"70",x"87"),
  1366 => (x"c0",x"87",x"d9",x"02"),
  1367 => (x"d3",x"02",x"ac",x"fb"),
  1368 => (x"ff",x"55",x"74",x"87"),
  1369 => (x"70",x"87",x"e1",x"dc"),
  1370 => (x"c7",x"02",x"9c",x"4c"),
  1371 => (x"ac",x"fb",x"c0",x"87"),
  1372 => (x"87",x"ed",x"ff",x"05"),
  1373 => (x"c2",x"55",x"e0",x"c0"),
  1374 => (x"97",x"c0",x"55",x"c1"),
  1375 => (x"66",x"e0",x"c0",x"7d"),
  1376 => (x"a8",x"66",x"c4",x"48"),
  1377 => (x"d0",x"87",x"db",x"05"),
  1378 => (x"66",x"d4",x"48",x"66"),
  1379 => (x"87",x"ca",x"04",x"a8"),
  1380 => (x"c1",x"48",x"66",x"d0"),
  1381 => (x"58",x"a6",x"d4",x"80"),
  1382 => (x"66",x"d4",x"87",x"c8"),
  1383 => (x"d8",x"88",x"c1",x"48"),
  1384 => (x"db",x"ff",x"58",x"a6"),
  1385 => (x"4c",x"70",x"87",x"e2"),
  1386 => (x"05",x"ac",x"d0",x"c1"),
  1387 => (x"66",x"dc",x"87",x"c9"),
  1388 => (x"c0",x"80",x"c1",x"48"),
  1389 => (x"c1",x"58",x"a6",x"e0"),
  1390 => (x"fd",x"02",x"ac",x"d0"),
  1391 => (x"48",x"6e",x"87",x"d9"),
  1392 => (x"a8",x"66",x"e0",x"c0"),
  1393 => (x"87",x"eb",x"c9",x"05"),
  1394 => (x"48",x"a6",x"e4",x"c0"),
  1395 => (x"48",x"74",x"78",x"c0"),
  1396 => (x"c8",x"88",x"fb",x"c0"),
  1397 => (x"98",x"70",x"58",x"a6"),
  1398 => (x"87",x"dd",x"c9",x"02"),
  1399 => (x"c8",x"88",x"cb",x"48"),
  1400 => (x"98",x"70",x"58",x"a6"),
  1401 => (x"87",x"cf",x"c1",x"02"),
  1402 => (x"c8",x"88",x"c9",x"48"),
  1403 => (x"98",x"70",x"58",x"a6"),
  1404 => (x"87",x"ff",x"c3",x"02"),
  1405 => (x"c8",x"88",x"c4",x"48"),
  1406 => (x"98",x"70",x"58",x"a6"),
  1407 => (x"48",x"87",x"cf",x"02"),
  1408 => (x"a6",x"c8",x"88",x"c1"),
  1409 => (x"02",x"98",x"70",x"58"),
  1410 => (x"c8",x"87",x"e8",x"c3"),
  1411 => (x"a6",x"c8",x"87",x"dc"),
  1412 => (x"78",x"f0",x"c0",x"48"),
  1413 => (x"87",x"f0",x"d9",x"ff"),
  1414 => (x"ec",x"c0",x"4c",x"70"),
  1415 => (x"c3",x"c0",x"02",x"ac"),
  1416 => (x"5c",x"a6",x"cc",x"87"),
  1417 => (x"02",x"ac",x"ec",x"c0"),
  1418 => (x"d9",x"ff",x"87",x"cd"),
  1419 => (x"4c",x"70",x"87",x"da"),
  1420 => (x"05",x"ac",x"ec",x"c0"),
  1421 => (x"c0",x"87",x"f3",x"ff"),
  1422 => (x"c0",x"02",x"ac",x"ec"),
  1423 => (x"d9",x"ff",x"87",x"c4"),
  1424 => (x"1e",x"c0",x"87",x"c6"),
  1425 => (x"66",x"d8",x"1e",x"ca"),
  1426 => (x"c1",x"91",x"cc",x"49"),
  1427 => (x"71",x"48",x"66",x"cc"),
  1428 => (x"58",x"a6",x"cc",x"80"),
  1429 => (x"c4",x"48",x"66",x"c8"),
  1430 => (x"58",x"a6",x"d0",x"80"),
  1431 => (x"49",x"bf",x"66",x"cc"),
  1432 => (x"87",x"e0",x"d9",x"ff"),
  1433 => (x"1e",x"de",x"1e",x"c1"),
  1434 => (x"49",x"bf",x"66",x"d4"),
  1435 => (x"87",x"d4",x"d9",x"ff"),
  1436 => (x"49",x"70",x"86",x"d0"),
  1437 => (x"88",x"08",x"c0",x"48"),
  1438 => (x"58",x"a6",x"ec",x"c0"),
  1439 => (x"c0",x"06",x"a8",x"c0"),
  1440 => (x"e8",x"c0",x"87",x"ee"),
  1441 => (x"a8",x"dd",x"48",x"66"),
  1442 => (x"87",x"e4",x"c0",x"03"),
  1443 => (x"49",x"bf",x"66",x"c4"),
  1444 => (x"81",x"66",x"e8",x"c0"),
  1445 => (x"c0",x"51",x"e0",x"c0"),
  1446 => (x"c1",x"49",x"66",x"e8"),
  1447 => (x"bf",x"66",x"c4",x"81"),
  1448 => (x"51",x"c1",x"c2",x"81"),
  1449 => (x"49",x"66",x"e8",x"c0"),
  1450 => (x"66",x"c4",x"81",x"c2"),
  1451 => (x"51",x"c0",x"81",x"bf"),
  1452 => (x"cb",x"c1",x"48",x"6e"),
  1453 => (x"49",x"6e",x"78",x"ce"),
  1454 => (x"66",x"d8",x"81",x"c8"),
  1455 => (x"c9",x"49",x"6e",x"51"),
  1456 => (x"51",x"66",x"dc",x"81"),
  1457 => (x"81",x"ca",x"49",x"6e"),
  1458 => (x"d8",x"51",x"66",x"c8"),
  1459 => (x"80",x"c1",x"48",x"66"),
  1460 => (x"d0",x"58",x"a6",x"dc"),
  1461 => (x"66",x"d4",x"48",x"66"),
  1462 => (x"cb",x"c0",x"04",x"a8"),
  1463 => (x"48",x"66",x"d0",x"87"),
  1464 => (x"a6",x"d4",x"80",x"c1"),
  1465 => (x"87",x"d1",x"c5",x"58"),
  1466 => (x"c1",x"48",x"66",x"d4"),
  1467 => (x"58",x"a6",x"d8",x"88"),
  1468 => (x"ff",x"87",x"c6",x"c5"),
  1469 => (x"c0",x"87",x"f8",x"d8"),
  1470 => (x"ff",x"58",x"a6",x"ec"),
  1471 => (x"c0",x"87",x"f0",x"d8"),
  1472 => (x"c0",x"58",x"a6",x"f0"),
  1473 => (x"c0",x"05",x"a8",x"ec"),
  1474 => (x"48",x"a6",x"87",x"c9"),
  1475 => (x"78",x"66",x"e8",x"c0"),
  1476 => (x"ff",x"87",x"c4",x"c0"),
  1477 => (x"d0",x"87",x"f1",x"d5"),
  1478 => (x"91",x"cc",x"49",x"66"),
  1479 => (x"48",x"66",x"c4",x"c1"),
  1480 => (x"a6",x"c8",x"80",x"71"),
  1481 => (x"4a",x"66",x"c4",x"58"),
  1482 => (x"66",x"c4",x"82",x"c8"),
  1483 => (x"c0",x"81",x"ca",x"49"),
  1484 => (x"c0",x"51",x"66",x"e8"),
  1485 => (x"c1",x"49",x"66",x"ec"),
  1486 => (x"66",x"e8",x"c0",x"81"),
  1487 => (x"71",x"48",x"c1",x"89"),
  1488 => (x"c1",x"49",x"70",x"30"),
  1489 => (x"7a",x"97",x"71",x"89"),
  1490 => (x"bf",x"e8",x"e3",x"c2"),
  1491 => (x"66",x"e8",x"c0",x"49"),
  1492 => (x"4a",x"6a",x"97",x"29"),
  1493 => (x"c0",x"98",x"71",x"48"),
  1494 => (x"c4",x"58",x"a6",x"f4"),
  1495 => (x"80",x"c4",x"48",x"66"),
  1496 => (x"c8",x"58",x"a6",x"cc"),
  1497 => (x"c0",x"4d",x"bf",x"66"),
  1498 => (x"6e",x"48",x"66",x"e0"),
  1499 => (x"c5",x"c0",x"02",x"a8"),
  1500 => (x"c0",x"7e",x"c0",x"87"),
  1501 => (x"7e",x"c1",x"87",x"c2"),
  1502 => (x"e0",x"c0",x"1e",x"6e"),
  1503 => (x"ff",x"49",x"75",x"1e"),
  1504 => (x"c8",x"87",x"c1",x"d5"),
  1505 => (x"c0",x"4c",x"70",x"86"),
  1506 => (x"c1",x"06",x"ac",x"b7"),
  1507 => (x"85",x"74",x"87",x"d4"),
  1508 => (x"49",x"bf",x"66",x"c8"),
  1509 => (x"75",x"81",x"e0",x"c0"),
  1510 => (x"c1",x"c1",x"4b",x"89"),
  1511 => (x"fe",x"71",x"4a",x"e0"),
  1512 => (x"c2",x"87",x"c0",x"e6"),
  1513 => (x"c0",x"7e",x"75",x"85"),
  1514 => (x"c1",x"48",x"66",x"e4"),
  1515 => (x"a6",x"e8",x"c0",x"80"),
  1516 => (x"66",x"f0",x"c0",x"58"),
  1517 => (x"70",x"81",x"c1",x"49"),
  1518 => (x"c5",x"c0",x"02",x"a9"),
  1519 => (x"c0",x"4d",x"c0",x"87"),
  1520 => (x"4d",x"c1",x"87",x"c2"),
  1521 => (x"66",x"cc",x"1e",x"75"),
  1522 => (x"e0",x"c0",x"49",x"bf"),
  1523 => (x"89",x"66",x"c4",x"81"),
  1524 => (x"66",x"c8",x"1e",x"71"),
  1525 => (x"eb",x"d3",x"ff",x"49"),
  1526 => (x"c0",x"86",x"c8",x"87"),
  1527 => (x"ff",x"01",x"a8",x"b7"),
  1528 => (x"e4",x"c0",x"87",x"c5"),
  1529 => (x"d3",x"c0",x"02",x"66"),
  1530 => (x"49",x"66",x"c4",x"87"),
  1531 => (x"e4",x"c0",x"81",x"c9"),
  1532 => (x"66",x"c4",x"51",x"66"),
  1533 => (x"e2",x"cd",x"c1",x"48"),
  1534 => (x"87",x"ce",x"c0",x"78"),
  1535 => (x"c9",x"49",x"66",x"c4"),
  1536 => (x"c4",x"51",x"c2",x"81"),
  1537 => (x"cf",x"c1",x"48",x"66"),
  1538 => (x"66",x"d0",x"78",x"e0"),
  1539 => (x"a8",x"66",x"d4",x"48"),
  1540 => (x"87",x"cb",x"c0",x"04"),
  1541 => (x"c1",x"48",x"66",x"d0"),
  1542 => (x"58",x"a6",x"d4",x"80"),
  1543 => (x"d4",x"87",x"da",x"c0"),
  1544 => (x"88",x"c1",x"48",x"66"),
  1545 => (x"c0",x"58",x"a6",x"d8"),
  1546 => (x"d2",x"ff",x"87",x"cf"),
  1547 => (x"4c",x"70",x"87",x"c2"),
  1548 => (x"ff",x"87",x"c6",x"c0"),
  1549 => (x"70",x"87",x"f9",x"d1"),
  1550 => (x"48",x"66",x"dc",x"4c"),
  1551 => (x"e0",x"c0",x"80",x"c1"),
  1552 => (x"9c",x"74",x"58",x"a6"),
  1553 => (x"87",x"cb",x"c0",x"02"),
  1554 => (x"c1",x"48",x"66",x"d0"),
  1555 => (x"04",x"a8",x"66",x"cc"),
  1556 => (x"d0",x"87",x"f1",x"f2"),
  1557 => (x"a8",x"c7",x"48",x"66"),
  1558 => (x"87",x"e1",x"c0",x"03"),
  1559 => (x"c2",x"4c",x"66",x"d0"),
  1560 => (x"c0",x"48",x"cc",x"e4"),
  1561 => (x"cc",x"49",x"74",x"78"),
  1562 => (x"66",x"c4",x"c1",x"91"),
  1563 => (x"4a",x"a1",x"c4",x"81"),
  1564 => (x"52",x"c0",x"4a",x"6a"),
  1565 => (x"c7",x"84",x"c1",x"79"),
  1566 => (x"e2",x"ff",x"04",x"ac"),
  1567 => (x"66",x"e0",x"c0",x"87"),
  1568 => (x"87",x"e2",x"c0",x"02"),
  1569 => (x"49",x"66",x"c4",x"c1"),
  1570 => (x"c1",x"81",x"d4",x"c1"),
  1571 => (x"c1",x"4a",x"66",x"c4"),
  1572 => (x"52",x"c0",x"82",x"dc"),
  1573 => (x"79",x"d4",x"cc",x"c1"),
  1574 => (x"49",x"66",x"c4",x"c1"),
  1575 => (x"c1",x"81",x"d8",x"c1"),
  1576 => (x"c0",x"79",x"e4",x"c1"),
  1577 => (x"c4",x"c1",x"87",x"d6"),
  1578 => (x"d4",x"c1",x"49",x"66"),
  1579 => (x"66",x"c4",x"c1",x"81"),
  1580 => (x"82",x"d8",x"c1",x"4a"),
  1581 => (x"7a",x"ec",x"c1",x"c1"),
  1582 => (x"79",x"cb",x"cc",x"c1"),
  1583 => (x"49",x"66",x"c4",x"c1"),
  1584 => (x"c1",x"81",x"e0",x"c1"),
  1585 => (x"ff",x"79",x"f2",x"cf"),
  1586 => (x"cc",x"87",x"dc",x"cf"),
  1587 => (x"cc",x"ff",x"48",x"66"),
  1588 => (x"26",x"4d",x"26",x"8e"),
  1589 => (x"26",x"4b",x"26",x"4c"),
  1590 => (x"1e",x"c7",x"1e",x"4f"),
  1591 => (x"bf",x"c8",x"e4",x"c2"),
  1592 => (x"d0",x"e6",x"c1",x"1e"),
  1593 => (x"ec",x"e3",x"c2",x"1e"),
  1594 => (x"ed",x"49",x"bf",x"97"),
  1595 => (x"e6",x"c1",x"87",x"d6"),
  1596 => (x"e1",x"c0",x"49",x"d0"),
  1597 => (x"8e",x"f4",x"87",x"f0"),
  1598 => (x"c1",x"1e",x"4f",x"26"),
  1599 => (x"c0",x"48",x"c4",x"e6"),
  1600 => (x"f0",x"d5",x"c2",x"50"),
  1601 => (x"d4",x"ff",x"49",x"bf"),
  1602 => (x"48",x"c0",x"87",x"d4"),
  1603 => (x"73",x"1e",x"4f",x"26"),
  1604 => (x"87",x"d9",x"c7",x"1e"),
  1605 => (x"48",x"d4",x"e4",x"c2"),
  1606 => (x"d4",x"ff",x"50",x"c0"),
  1607 => (x"78",x"ff",x"c3",x"48"),
  1608 => (x"49",x"f4",x"c1",x"c1"),
  1609 => (x"87",x"ff",x"dd",x"fe"),
  1610 => (x"87",x"d4",x"e9",x"fe"),
  1611 => (x"cd",x"02",x"98",x"70"),
  1612 => (x"c7",x"f1",x"fe",x"87"),
  1613 => (x"02",x"98",x"70",x"87"),
  1614 => (x"4a",x"c1",x"87",x"c4"),
  1615 => (x"4a",x"c0",x"87",x"c2"),
  1616 => (x"c8",x"02",x"9a",x"72"),
  1617 => (x"c0",x"c2",x"c1",x"87"),
  1618 => (x"da",x"dd",x"fe",x"49"),
  1619 => (x"c8",x"e4",x"c2",x"87"),
  1620 => (x"c2",x"78",x"c0",x"48"),
  1621 => (x"c0",x"48",x"ec",x"e3"),
  1622 => (x"fc",x"fd",x"49",x"50"),
  1623 => (x"87",x"da",x"fe",x"87"),
  1624 => (x"02",x"9b",x"4b",x"70"),
  1625 => (x"e7",x"c1",x"87",x"cf"),
  1626 => (x"49",x"c7",x"5b",x"ec"),
  1627 => (x"c1",x"87",x"e9",x"de"),
  1628 => (x"c4",x"e0",x"c0",x"49"),
  1629 => (x"87",x"ef",x"c2",x"87"),
  1630 => (x"87",x"e5",x"e1",x"c0"),
  1631 => (x"4b",x"26",x"87",x"fa"),
  1632 => (x"00",x"00",x"4f",x"26"),
  1633 => (x"00",x"00",x"00",x"00"),
  1634 => (x"00",x"00",x"00",x"00"),
  1635 => (x"00",x"00",x"00",x"01"),
  1636 => (x"00",x"00",x"0f",x"be"),
  1637 => (x"00",x"00",x"29",x"20"),
  1638 => (x"00",x"00",x"00",x"00"),
  1639 => (x"00",x"00",x"0f",x"be"),
  1640 => (x"00",x"00",x"29",x"3e"),
  1641 => (x"00",x"00",x"00",x"00"),
  1642 => (x"00",x"00",x"0f",x"be"),
  1643 => (x"00",x"00",x"29",x"5c"),
  1644 => (x"00",x"00",x"00",x"00"),
  1645 => (x"00",x"00",x"0f",x"be"),
  1646 => (x"00",x"00",x"29",x"7a"),
  1647 => (x"00",x"00",x"00",x"00"),
  1648 => (x"00",x"00",x"0f",x"be"),
  1649 => (x"00",x"00",x"29",x"98"),
  1650 => (x"00",x"00",x"00",x"00"),
  1651 => (x"00",x"00",x"0f",x"be"),
  1652 => (x"00",x"00",x"29",x"b6"),
  1653 => (x"00",x"00",x"00",x"00"),
  1654 => (x"00",x"00",x"0f",x"be"),
  1655 => (x"00",x"00",x"29",x"d4"),
  1656 => (x"00",x"00",x"00",x"00"),
  1657 => (x"00",x"00",x"13",x"14"),
  1658 => (x"00",x"00",x"00",x"00"),
  1659 => (x"00",x"00",x"00",x"00"),
  1660 => (x"00",x"00",x"10",x"b8"),
  1661 => (x"00",x"00",x"00",x"00"),
  1662 => (x"00",x"00",x"00",x"00"),
  1663 => (x"00",x"00",x"10",x"84"),
  1664 => (x"db",x"86",x"fc",x"1e"),
  1665 => (x"fc",x"7e",x"70",x"87"),
  1666 => (x"1e",x"4f",x"26",x"8e"),
  1667 => (x"c0",x"48",x"f0",x"fe"),
  1668 => (x"79",x"09",x"cd",x"78"),
  1669 => (x"1e",x"4f",x"26",x"09"),
  1670 => (x"49",x"c0",x"e8",x"c1"),
  1671 => (x"4f",x"26",x"87",x"ed"),
  1672 => (x"bf",x"f0",x"fe",x"1e"),
  1673 => (x"1e",x"4f",x"26",x"48"),
  1674 => (x"c1",x"48",x"f0",x"fe"),
  1675 => (x"1e",x"4f",x"26",x"78"),
  1676 => (x"c0",x"48",x"f0",x"fe"),
  1677 => (x"1e",x"4f",x"26",x"78"),
  1678 => (x"52",x"c0",x"4a",x"71"),
  1679 => (x"0e",x"4f",x"26",x"51"),
  1680 => (x"5d",x"5c",x"5b",x"5e"),
  1681 => (x"71",x"86",x"f4",x"0e"),
  1682 => (x"7e",x"6d",x"97",x"4d"),
  1683 => (x"97",x"4c",x"a5",x"c1"),
  1684 => (x"a6",x"c8",x"48",x"6c"),
  1685 => (x"c4",x"48",x"6e",x"58"),
  1686 => (x"c5",x"05",x"a8",x"66"),
  1687 => (x"c0",x"48",x"ff",x"87"),
  1688 => (x"ca",x"ff",x"87",x"e6"),
  1689 => (x"49",x"a5",x"c2",x"87"),
  1690 => (x"71",x"4b",x"6c",x"97"),
  1691 => (x"6b",x"97",x"4b",x"a3"),
  1692 => (x"7e",x"6c",x"97",x"4b"),
  1693 => (x"80",x"c1",x"48",x"6e"),
  1694 => (x"c7",x"58",x"a6",x"c8"),
  1695 => (x"58",x"a6",x"cc",x"98"),
  1696 => (x"fe",x"7c",x"97",x"70"),
  1697 => (x"48",x"73",x"87",x"e1"),
  1698 => (x"4d",x"26",x"8e",x"f4"),
  1699 => (x"4b",x"26",x"4c",x"26"),
  1700 => (x"5e",x"0e",x"4f",x"26"),
  1701 => (x"f4",x"0e",x"5c",x"5b"),
  1702 => (x"d8",x"4c",x"71",x"86"),
  1703 => (x"ff",x"c3",x"4a",x"66"),
  1704 => (x"4b",x"a4",x"c2",x"9a"),
  1705 => (x"73",x"49",x"6c",x"97"),
  1706 => (x"51",x"72",x"49",x"a1"),
  1707 => (x"6e",x"7e",x"6c",x"97"),
  1708 => (x"c8",x"80",x"c1",x"48"),
  1709 => (x"98",x"c7",x"58",x"a6"),
  1710 => (x"70",x"58",x"a6",x"cc"),
  1711 => (x"26",x"8e",x"f4",x"54"),
  1712 => (x"26",x"4b",x"26",x"4c"),
  1713 => (x"86",x"fc",x"1e",x"4f"),
  1714 => (x"e0",x"87",x"e4",x"fd"),
  1715 => (x"c0",x"49",x"4a",x"bf"),
  1716 => (x"02",x"99",x"c0",x"e0"),
  1717 => (x"1e",x"72",x"87",x"cb"),
  1718 => (x"49",x"c8",x"e8",x"c2"),
  1719 => (x"c4",x"87",x"f3",x"fe"),
  1720 => (x"87",x"fc",x"fc",x"86"),
  1721 => (x"fe",x"fc",x"7e",x"70"),
  1722 => (x"26",x"8e",x"fc",x"87"),
  1723 => (x"e8",x"c2",x"1e",x"4f"),
  1724 => (x"c2",x"fd",x"49",x"c8"),
  1725 => (x"c5",x"eb",x"c1",x"87"),
  1726 => (x"87",x"cf",x"fc",x"49"),
  1727 => (x"26",x"87",x"ed",x"c4"),
  1728 => (x"5b",x"5e",x"0e",x"4f"),
  1729 => (x"fc",x"0e",x"5d",x"5c"),
  1730 => (x"ff",x"7e",x"71",x"86"),
  1731 => (x"e8",x"c2",x"4d",x"d4"),
  1732 => (x"ea",x"fc",x"49",x"c8"),
  1733 => (x"c0",x"4b",x"70",x"87"),
  1734 => (x"c2",x"04",x"ab",x"b7"),
  1735 => (x"f0",x"c3",x"87",x"f8"),
  1736 => (x"87",x"c9",x"05",x"ab"),
  1737 => (x"48",x"e4",x"ef",x"c1"),
  1738 => (x"d9",x"c2",x"78",x"c1"),
  1739 => (x"ab",x"e0",x"c3",x"87"),
  1740 => (x"c1",x"87",x"c9",x"05"),
  1741 => (x"c1",x"48",x"e8",x"ef"),
  1742 => (x"87",x"ca",x"c2",x"78"),
  1743 => (x"bf",x"e8",x"ef",x"c1"),
  1744 => (x"c2",x"87",x"c6",x"02"),
  1745 => (x"c2",x"4c",x"a3",x"c0"),
  1746 => (x"c1",x"4c",x"73",x"87"),
  1747 => (x"02",x"bf",x"e4",x"ef"),
  1748 => (x"74",x"87",x"e0",x"c0"),
  1749 => (x"29",x"b7",x"c4",x"49"),
  1750 => (x"ec",x"ef",x"c1",x"91"),
  1751 => (x"cf",x"4a",x"74",x"81"),
  1752 => (x"c1",x"92",x"c2",x"9a"),
  1753 => (x"70",x"30",x"72",x"48"),
  1754 => (x"72",x"ba",x"ff",x"4a"),
  1755 => (x"70",x"98",x"69",x"48"),
  1756 => (x"74",x"87",x"db",x"79"),
  1757 => (x"29",x"b7",x"c4",x"49"),
  1758 => (x"ec",x"ef",x"c1",x"91"),
  1759 => (x"cf",x"4a",x"74",x"81"),
  1760 => (x"c3",x"92",x"c2",x"9a"),
  1761 => (x"70",x"30",x"72",x"48"),
  1762 => (x"b0",x"69",x"48",x"4a"),
  1763 => (x"05",x"6e",x"79",x"70"),
  1764 => (x"ff",x"87",x"e7",x"c0"),
  1765 => (x"e1",x"c8",x"48",x"d0"),
  1766 => (x"c1",x"7d",x"c5",x"78"),
  1767 => (x"02",x"bf",x"e8",x"ef"),
  1768 => (x"e0",x"c3",x"87",x"c3"),
  1769 => (x"e4",x"ef",x"c1",x"7d"),
  1770 => (x"87",x"c3",x"02",x"bf"),
  1771 => (x"73",x"7d",x"f0",x"c3"),
  1772 => (x"48",x"d0",x"ff",x"7d"),
  1773 => (x"c0",x"78",x"e1",x"c8"),
  1774 => (x"ef",x"c1",x"78",x"e0"),
  1775 => (x"78",x"c0",x"48",x"e8"),
  1776 => (x"48",x"e4",x"ef",x"c1"),
  1777 => (x"e8",x"c2",x"78",x"c0"),
  1778 => (x"f2",x"f9",x"49",x"c8"),
  1779 => (x"c0",x"4b",x"70",x"87"),
  1780 => (x"fd",x"03",x"ab",x"b7"),
  1781 => (x"48",x"c0",x"87",x"c8"),
  1782 => (x"4d",x"26",x"8e",x"fc"),
  1783 => (x"4b",x"26",x"4c",x"26"),
  1784 => (x"00",x"00",x"4f",x"26"),
  1785 => (x"00",x"00",x"00",x"00"),
  1786 => (x"00",x"00",x"00",x"00"),
  1787 => (x"00",x"00",x"00",x"00"),
  1788 => (x"00",x"00",x"00",x"00"),
  1789 => (x"00",x"00",x"00",x"00"),
  1790 => (x"00",x"00",x"00",x"00"),
  1791 => (x"00",x"00",x"00",x"00"),
  1792 => (x"00",x"00",x"00",x"00"),
  1793 => (x"00",x"00",x"00",x"00"),
  1794 => (x"00",x"00",x"00",x"00"),
  1795 => (x"00",x"00",x"00",x"00"),
  1796 => (x"00",x"00",x"00",x"00"),
  1797 => (x"00",x"00",x"00",x"00"),
  1798 => (x"00",x"00",x"00",x"00"),
  1799 => (x"00",x"00",x"00",x"00"),
  1800 => (x"00",x"00",x"00",x"00"),
  1801 => (x"00",x"00",x"00",x"00"),
  1802 => (x"00",x"00",x"00",x"00"),
  1803 => (x"72",x"4a",x"c0",x"1e"),
  1804 => (x"c1",x"91",x"c4",x"49"),
  1805 => (x"c0",x"81",x"ec",x"ef"),
  1806 => (x"d0",x"82",x"c1",x"79"),
  1807 => (x"ee",x"04",x"aa",x"b7"),
  1808 => (x"0e",x"4f",x"26",x"87"),
  1809 => (x"5d",x"5c",x"5b",x"5e"),
  1810 => (x"f7",x"4d",x"71",x"0e"),
  1811 => (x"4a",x"75",x"87",x"e1"),
  1812 => (x"92",x"2a",x"b7",x"c4"),
  1813 => (x"82",x"ec",x"ef",x"c1"),
  1814 => (x"9c",x"cf",x"4c",x"75"),
  1815 => (x"49",x"6a",x"94",x"c2"),
  1816 => (x"c3",x"2b",x"74",x"4b"),
  1817 => (x"74",x"48",x"c2",x"9b"),
  1818 => (x"ff",x"4c",x"70",x"30"),
  1819 => (x"71",x"48",x"74",x"bc"),
  1820 => (x"f6",x"7a",x"70",x"98"),
  1821 => (x"48",x"73",x"87",x"f1"),
  1822 => (x"4c",x"26",x"4d",x"26"),
  1823 => (x"4f",x"26",x"4b",x"26"),
  1824 => (x"48",x"d0",x"ff",x"1e"),
  1825 => (x"71",x"78",x"e1",x"c8"),
  1826 => (x"08",x"d4",x"ff",x"48"),
  1827 => (x"48",x"66",x"c4",x"78"),
  1828 => (x"78",x"08",x"d4",x"ff"),
  1829 => (x"71",x"1e",x"4f",x"26"),
  1830 => (x"49",x"66",x"c4",x"4a"),
  1831 => (x"ff",x"49",x"72",x"1e"),
  1832 => (x"d0",x"ff",x"87",x"de"),
  1833 => (x"78",x"e0",x"c0",x"48"),
  1834 => (x"4f",x"26",x"8e",x"fc"),
  1835 => (x"71",x"1e",x"73",x"1e"),
  1836 => (x"49",x"66",x"c8",x"4b"),
  1837 => (x"c1",x"4a",x"73",x"1e"),
  1838 => (x"ff",x"49",x"a2",x"e0"),
  1839 => (x"8e",x"fc",x"87",x"d8"),
  1840 => (x"4f",x"26",x"4b",x"26"),
  1841 => (x"48",x"d0",x"ff",x"1e"),
  1842 => (x"71",x"78",x"c9",x"c8"),
  1843 => (x"08",x"d4",x"ff",x"48"),
  1844 => (x"1e",x"4f",x"26",x"78"),
  1845 => (x"eb",x"49",x"4a",x"71"),
  1846 => (x"48",x"d0",x"ff",x"87"),
  1847 => (x"4f",x"26",x"78",x"c8"),
  1848 => (x"71",x"1e",x"73",x"1e"),
  1849 => (x"e0",x"e8",x"c2",x"4b"),
  1850 => (x"87",x"c3",x"02",x"bf"),
  1851 => (x"ff",x"87",x"eb",x"c2"),
  1852 => (x"c9",x"c8",x"48",x"d0"),
  1853 => (x"c0",x"48",x"73",x"78"),
  1854 => (x"d4",x"ff",x"b0",x"e0"),
  1855 => (x"e8",x"c2",x"78",x"08"),
  1856 => (x"78",x"c0",x"48",x"d4"),
  1857 => (x"c5",x"02",x"66",x"c8"),
  1858 => (x"49",x"ff",x"c3",x"87"),
  1859 => (x"49",x"c0",x"87",x"c2"),
  1860 => (x"59",x"dc",x"e8",x"c2"),
  1861 => (x"c6",x"02",x"66",x"cc"),
  1862 => (x"d5",x"d5",x"c5",x"87"),
  1863 => (x"cf",x"87",x"c4",x"4a"),
  1864 => (x"c2",x"4a",x"ff",x"ff"),
  1865 => (x"c2",x"5a",x"e0",x"e8"),
  1866 => (x"c1",x"48",x"e0",x"e8"),
  1867 => (x"26",x"4b",x"26",x"78"),
  1868 => (x"5b",x"5e",x"0e",x"4f"),
  1869 => (x"71",x"0e",x"5d",x"5c"),
  1870 => (x"dc",x"e8",x"c2",x"4d"),
  1871 => (x"9d",x"75",x"4b",x"bf"),
  1872 => (x"49",x"87",x"cb",x"02"),
  1873 => (x"f3",x"c1",x"91",x"c8"),
  1874 => (x"82",x"71",x"4a",x"d8"),
  1875 => (x"f7",x"c1",x"87",x"c4"),
  1876 => (x"4c",x"c0",x"4a",x"d8"),
  1877 => (x"99",x"73",x"49",x"12"),
  1878 => (x"bf",x"d8",x"e8",x"c2"),
  1879 => (x"ff",x"b8",x"71",x"48"),
  1880 => (x"c1",x"78",x"08",x"d4"),
  1881 => (x"c8",x"84",x"2b",x"b7"),
  1882 => (x"e7",x"04",x"ac",x"b7"),
  1883 => (x"d4",x"e8",x"c2",x"87"),
  1884 => (x"80",x"c8",x"48",x"bf"),
  1885 => (x"58",x"d8",x"e8",x"c2"),
  1886 => (x"4c",x"26",x"4d",x"26"),
  1887 => (x"4f",x"26",x"4b",x"26"),
  1888 => (x"71",x"1e",x"73",x"1e"),
  1889 => (x"9a",x"4a",x"13",x"4b"),
  1890 => (x"72",x"87",x"cb",x"02"),
  1891 => (x"87",x"e1",x"fe",x"49"),
  1892 => (x"05",x"9a",x"4a",x"13"),
  1893 => (x"4b",x"26",x"87",x"f5"),
  1894 => (x"c2",x"1e",x"4f",x"26"),
  1895 => (x"49",x"bf",x"d4",x"e8"),
  1896 => (x"48",x"d4",x"e8",x"c2"),
  1897 => (x"c4",x"78",x"a1",x"c1"),
  1898 => (x"03",x"a9",x"b7",x"c0"),
  1899 => (x"d4",x"ff",x"87",x"db"),
  1900 => (x"d8",x"e8",x"c2",x"48"),
  1901 => (x"e8",x"c2",x"78",x"bf"),
  1902 => (x"c2",x"49",x"bf",x"d4"),
  1903 => (x"c1",x"48",x"d4",x"e8"),
  1904 => (x"c0",x"c4",x"78",x"a1"),
  1905 => (x"e5",x"04",x"a9",x"b7"),
  1906 => (x"48",x"d0",x"ff",x"87"),
  1907 => (x"e8",x"c2",x"78",x"c8"),
  1908 => (x"78",x"c0",x"48",x"e0"),
  1909 => (x"00",x"00",x"4f",x"26"),
  1910 => (x"00",x"00",x"00",x"00"),
  1911 => (x"00",x"00",x"00",x"00"),
  1912 => (x"5f",x"00",x"00",x"00"),
  1913 => (x"00",x"00",x"00",x"5f"),
  1914 => (x"00",x"03",x"03",x"00"),
  1915 => (x"00",x"00",x"03",x"03"),
  1916 => (x"14",x"7f",x"7f",x"14"),
  1917 => (x"00",x"14",x"7f",x"7f"),
  1918 => (x"6b",x"2e",x"24",x"00"),
  1919 => (x"00",x"12",x"3a",x"6b"),
  1920 => (x"18",x"36",x"6a",x"4c"),
  1921 => (x"00",x"32",x"56",x"6c"),
  1922 => (x"59",x"4f",x"7e",x"30"),
  1923 => (x"40",x"68",x"3a",x"77"),
  1924 => (x"07",x"04",x"00",x"00"),
  1925 => (x"00",x"00",x"00",x"03"),
  1926 => (x"3e",x"1c",x"00",x"00"),
  1927 => (x"00",x"00",x"41",x"63"),
  1928 => (x"63",x"41",x"00",x"00"),
  1929 => (x"00",x"00",x"1c",x"3e"),
  1930 => (x"1c",x"3e",x"2a",x"08"),
  1931 => (x"08",x"2a",x"3e",x"1c"),
  1932 => (x"3e",x"08",x"08",x"00"),
  1933 => (x"00",x"08",x"08",x"3e"),
  1934 => (x"e0",x"80",x"00",x"00"),
  1935 => (x"00",x"00",x"00",x"60"),
  1936 => (x"08",x"08",x"08",x"00"),
  1937 => (x"00",x"08",x"08",x"08"),
  1938 => (x"60",x"00",x"00",x"00"),
  1939 => (x"00",x"00",x"00",x"60"),
  1940 => (x"18",x"30",x"60",x"40"),
  1941 => (x"01",x"03",x"06",x"0c"),
  1942 => (x"59",x"7f",x"3e",x"00"),
  1943 => (x"00",x"3e",x"7f",x"4d"),
  1944 => (x"7f",x"06",x"04",x"00"),
  1945 => (x"00",x"00",x"00",x"7f"),
  1946 => (x"71",x"63",x"42",x"00"),
  1947 => (x"00",x"46",x"4f",x"59"),
  1948 => (x"49",x"63",x"22",x"00"),
  1949 => (x"00",x"36",x"7f",x"49"),
  1950 => (x"13",x"16",x"1c",x"18"),
  1951 => (x"00",x"10",x"7f",x"7f"),
  1952 => (x"45",x"67",x"27",x"00"),
  1953 => (x"00",x"39",x"7d",x"45"),
  1954 => (x"4b",x"7e",x"3c",x"00"),
  1955 => (x"00",x"30",x"79",x"49"),
  1956 => (x"71",x"01",x"01",x"00"),
  1957 => (x"00",x"07",x"0f",x"79"),
  1958 => (x"49",x"7f",x"36",x"00"),
  1959 => (x"00",x"36",x"7f",x"49"),
  1960 => (x"49",x"4f",x"06",x"00"),
  1961 => (x"00",x"1e",x"3f",x"69"),
  1962 => (x"66",x"00",x"00",x"00"),
  1963 => (x"00",x"00",x"00",x"66"),
  1964 => (x"e6",x"80",x"00",x"00"),
  1965 => (x"00",x"00",x"00",x"66"),
  1966 => (x"14",x"08",x"08",x"00"),
  1967 => (x"00",x"22",x"22",x"14"),
  1968 => (x"14",x"14",x"14",x"00"),
  1969 => (x"00",x"14",x"14",x"14"),
  1970 => (x"14",x"22",x"22",x"00"),
  1971 => (x"00",x"08",x"08",x"14"),
  1972 => (x"51",x"03",x"02",x"00"),
  1973 => (x"00",x"06",x"0f",x"59"),
  1974 => (x"5d",x"41",x"7f",x"3e"),
  1975 => (x"00",x"1e",x"1f",x"55"),
  1976 => (x"09",x"7f",x"7e",x"00"),
  1977 => (x"00",x"7e",x"7f",x"09"),
  1978 => (x"49",x"7f",x"7f",x"00"),
  1979 => (x"00",x"36",x"7f",x"49"),
  1980 => (x"63",x"3e",x"1c",x"00"),
  1981 => (x"00",x"41",x"41",x"41"),
  1982 => (x"41",x"7f",x"7f",x"00"),
  1983 => (x"00",x"1c",x"3e",x"63"),
  1984 => (x"49",x"7f",x"7f",x"00"),
  1985 => (x"00",x"41",x"41",x"49"),
  1986 => (x"09",x"7f",x"7f",x"00"),
  1987 => (x"00",x"01",x"01",x"09"),
  1988 => (x"41",x"7f",x"3e",x"00"),
  1989 => (x"00",x"7a",x"7b",x"49"),
  1990 => (x"08",x"7f",x"7f",x"00"),
  1991 => (x"00",x"7f",x"7f",x"08"),
  1992 => (x"7f",x"41",x"00",x"00"),
  1993 => (x"00",x"00",x"41",x"7f"),
  1994 => (x"40",x"60",x"20",x"00"),
  1995 => (x"00",x"3f",x"7f",x"40"),
  1996 => (x"1c",x"08",x"7f",x"7f"),
  1997 => (x"00",x"41",x"63",x"36"),
  1998 => (x"40",x"7f",x"7f",x"00"),
  1999 => (x"00",x"40",x"40",x"40"),
  2000 => (x"0c",x"06",x"7f",x"7f"),
  2001 => (x"00",x"7f",x"7f",x"06"),
  2002 => (x"0c",x"06",x"7f",x"7f"),
  2003 => (x"00",x"7f",x"7f",x"18"),
  2004 => (x"41",x"7f",x"3e",x"00"),
  2005 => (x"00",x"3e",x"7f",x"41"),
  2006 => (x"09",x"7f",x"7f",x"00"),
  2007 => (x"00",x"06",x"0f",x"09"),
  2008 => (x"61",x"41",x"7f",x"3e"),
  2009 => (x"00",x"40",x"7e",x"7f"),
  2010 => (x"09",x"7f",x"7f",x"00"),
  2011 => (x"00",x"66",x"7f",x"19"),
  2012 => (x"4d",x"6f",x"26",x"00"),
  2013 => (x"00",x"32",x"7b",x"59"),
  2014 => (x"7f",x"01",x"01",x"00"),
  2015 => (x"00",x"01",x"01",x"7f"),
  2016 => (x"40",x"7f",x"3f",x"00"),
  2017 => (x"00",x"3f",x"7f",x"40"),
  2018 => (x"70",x"3f",x"0f",x"00"),
  2019 => (x"00",x"0f",x"3f",x"70"),
  2020 => (x"18",x"30",x"7f",x"7f"),
  2021 => (x"00",x"7f",x"7f",x"30"),
  2022 => (x"1c",x"36",x"63",x"41"),
  2023 => (x"41",x"63",x"36",x"1c"),
  2024 => (x"7c",x"06",x"03",x"01"),
  2025 => (x"01",x"03",x"06",x"7c"),
  2026 => (x"4d",x"59",x"71",x"61"),
  2027 => (x"00",x"41",x"43",x"47"),
  2028 => (x"7f",x"7f",x"00",x"00"),
  2029 => (x"00",x"00",x"41",x"41"),
  2030 => (x"0c",x"06",x"03",x"01"),
  2031 => (x"40",x"60",x"30",x"18"),
  2032 => (x"41",x"41",x"00",x"00"),
  2033 => (x"00",x"00",x"7f",x"7f"),
  2034 => (x"03",x"06",x"0c",x"08"),
  2035 => (x"00",x"08",x"0c",x"06"),
  2036 => (x"80",x"80",x"80",x"80"),
  2037 => (x"00",x"80",x"80",x"80"),
  2038 => (x"03",x"00",x"00",x"00"),
  2039 => (x"00",x"00",x"04",x"07"),
  2040 => (x"54",x"74",x"20",x"00"),
  2041 => (x"00",x"78",x"7c",x"54"),
  2042 => (x"44",x"7f",x"7f",x"00"),
  2043 => (x"00",x"38",x"7c",x"44"),
  2044 => (x"44",x"7c",x"38",x"00"),
  2045 => (x"00",x"00",x"44",x"44"),
  2046 => (x"44",x"7c",x"38",x"00"),
  2047 => (x"00",x"7f",x"7f",x"44"),
  2048 => (x"54",x"7c",x"38",x"00"),
  2049 => (x"00",x"18",x"5c",x"54"),
  2050 => (x"7f",x"7e",x"04",x"00"),
  2051 => (x"00",x"00",x"05",x"05"),
  2052 => (x"a4",x"bc",x"18",x"00"),
  2053 => (x"00",x"7c",x"fc",x"a4"),
  2054 => (x"04",x"7f",x"7f",x"00"),
  2055 => (x"00",x"78",x"7c",x"04"),
  2056 => (x"3d",x"00",x"00",x"00"),
  2057 => (x"00",x"00",x"40",x"7d"),
  2058 => (x"80",x"80",x"80",x"00"),
  2059 => (x"00",x"00",x"7d",x"fd"),
  2060 => (x"10",x"7f",x"7f",x"00"),
  2061 => (x"00",x"44",x"6c",x"38"),
  2062 => (x"3f",x"00",x"00",x"00"),
  2063 => (x"00",x"00",x"40",x"7f"),
  2064 => (x"18",x"0c",x"7c",x"7c"),
  2065 => (x"00",x"78",x"7c",x"0c"),
  2066 => (x"04",x"7c",x"7c",x"00"),
  2067 => (x"00",x"78",x"7c",x"04"),
  2068 => (x"44",x"7c",x"38",x"00"),
  2069 => (x"00",x"38",x"7c",x"44"),
  2070 => (x"24",x"fc",x"fc",x"00"),
  2071 => (x"00",x"18",x"3c",x"24"),
  2072 => (x"24",x"3c",x"18",x"00"),
  2073 => (x"00",x"fc",x"fc",x"24"),
  2074 => (x"04",x"7c",x"7c",x"00"),
  2075 => (x"00",x"08",x"0c",x"04"),
  2076 => (x"54",x"5c",x"48",x"00"),
  2077 => (x"00",x"20",x"74",x"54"),
  2078 => (x"7f",x"3f",x"04",x"00"),
  2079 => (x"00",x"00",x"44",x"44"),
  2080 => (x"40",x"7c",x"3c",x"00"),
  2081 => (x"00",x"7c",x"7c",x"40"),
  2082 => (x"60",x"3c",x"1c",x"00"),
  2083 => (x"00",x"1c",x"3c",x"60"),
  2084 => (x"30",x"60",x"7c",x"3c"),
  2085 => (x"00",x"3c",x"7c",x"60"),
  2086 => (x"10",x"38",x"6c",x"44"),
  2087 => (x"00",x"44",x"6c",x"38"),
  2088 => (x"e0",x"bc",x"1c",x"00"),
  2089 => (x"00",x"1c",x"3c",x"60"),
  2090 => (x"74",x"64",x"44",x"00"),
  2091 => (x"00",x"44",x"4c",x"5c"),
  2092 => (x"3e",x"08",x"08",x"00"),
  2093 => (x"00",x"41",x"41",x"77"),
  2094 => (x"7f",x"00",x"00",x"00"),
  2095 => (x"00",x"00",x"00",x"7f"),
  2096 => (x"77",x"41",x"41",x"00"),
  2097 => (x"00",x"08",x"08",x"3e"),
  2098 => (x"03",x"01",x"01",x"02"),
  2099 => (x"00",x"01",x"02",x"02"),
  2100 => (x"7f",x"7f",x"7f",x"7f"),
  2101 => (x"00",x"7f",x"7f",x"7f"),
  2102 => (x"1c",x"1c",x"08",x"08"),
  2103 => (x"7f",x"7f",x"3e",x"3e"),
  2104 => (x"3e",x"3e",x"7f",x"7f"),
  2105 => (x"08",x"08",x"1c",x"1c"),
  2106 => (x"7c",x"18",x"10",x"00"),
  2107 => (x"00",x"10",x"18",x"7c"),
  2108 => (x"7c",x"30",x"10",x"00"),
  2109 => (x"00",x"10",x"30",x"7c"),
  2110 => (x"60",x"60",x"30",x"10"),
  2111 => (x"00",x"06",x"1e",x"78"),
  2112 => (x"18",x"3c",x"66",x"42"),
  2113 => (x"00",x"42",x"66",x"3c"),
  2114 => (x"c2",x"6a",x"38",x"78"),
  2115 => (x"00",x"38",x"6c",x"c6"),
  2116 => (x"60",x"00",x"00",x"60"),
  2117 => (x"00",x"60",x"00",x"00"),
  2118 => (x"5c",x"5b",x"5e",x"0e"),
  2119 => (x"86",x"fc",x"0e",x"5d"),
  2120 => (x"e8",x"c2",x"7e",x"71"),
  2121 => (x"c0",x"4c",x"bf",x"e8"),
  2122 => (x"c4",x"1e",x"c0",x"4b"),
  2123 => (x"c4",x"02",x"ab",x"66"),
  2124 => (x"c2",x"4d",x"c0",x"87"),
  2125 => (x"75",x"4d",x"c1",x"87"),
  2126 => (x"ee",x"49",x"73",x"1e"),
  2127 => (x"86",x"c8",x"87",x"e2"),
  2128 => (x"ef",x"49",x"e0",x"c0"),
  2129 => (x"a4",x"c4",x"87",x"eb"),
  2130 => (x"f0",x"49",x"6a",x"4a"),
  2131 => (x"c9",x"f1",x"87",x"f2"),
  2132 => (x"c1",x"84",x"cc",x"87"),
  2133 => (x"ab",x"b7",x"c8",x"83"),
  2134 => (x"87",x"cd",x"ff",x"04"),
  2135 => (x"4d",x"26",x"8e",x"fc"),
  2136 => (x"4b",x"26",x"4c",x"26"),
  2137 => (x"71",x"1e",x"4f",x"26"),
  2138 => (x"ec",x"e8",x"c2",x"4a"),
  2139 => (x"ec",x"e8",x"c2",x"5a"),
  2140 => (x"49",x"78",x"c7",x"48"),
  2141 => (x"26",x"87",x"e1",x"fe"),
  2142 => (x"1e",x"73",x"1e",x"4f"),
  2143 => (x"b7",x"c0",x"4a",x"71"),
  2144 => (x"87",x"d3",x"03",x"aa"),
  2145 => (x"bf",x"f4",x"d4",x"c2"),
  2146 => (x"c1",x"87",x"c4",x"05"),
  2147 => (x"c0",x"87",x"c2",x"4b"),
  2148 => (x"f8",x"d4",x"c2",x"4b"),
  2149 => (x"c2",x"87",x"c4",x"5b"),
  2150 => (x"fc",x"5a",x"f8",x"d4"),
  2151 => (x"f4",x"d4",x"c2",x"48"),
  2152 => (x"c1",x"4a",x"78",x"bf"),
  2153 => (x"a2",x"c0",x"c1",x"9a"),
  2154 => (x"87",x"e7",x"ec",x"49"),
  2155 => (x"4f",x"26",x"4b",x"26"),
  2156 => (x"c4",x"4a",x"71",x"1e"),
  2157 => (x"49",x"72",x"1e",x"66"),
  2158 => (x"fc",x"87",x"f1",x"eb"),
  2159 => (x"1e",x"4f",x"26",x"8e"),
  2160 => (x"c3",x"48",x"d4",x"ff"),
  2161 => (x"d0",x"ff",x"78",x"ff"),
  2162 => (x"78",x"e1",x"c0",x"48"),
  2163 => (x"c1",x"48",x"d4",x"ff"),
  2164 => (x"c4",x"48",x"71",x"78"),
  2165 => (x"08",x"d4",x"ff",x"30"),
  2166 => (x"48",x"d0",x"ff",x"78"),
  2167 => (x"26",x"78",x"e0",x"c0"),
  2168 => (x"5b",x"5e",x"0e",x"4f"),
  2169 => (x"f0",x"0e",x"5d",x"5c"),
  2170 => (x"48",x"a6",x"c8",x"86"),
  2171 => (x"bf",x"ec",x"78",x"c0"),
  2172 => (x"c2",x"80",x"fc",x"7e"),
  2173 => (x"78",x"bf",x"e8",x"e8"),
  2174 => (x"bf",x"f0",x"e8",x"c2"),
  2175 => (x"4c",x"bf",x"e8",x"4d"),
  2176 => (x"bf",x"f4",x"d4",x"c2"),
  2177 => (x"87",x"f9",x"e3",x"49"),
  2178 => (x"f6",x"e8",x"49",x"c7"),
  2179 => (x"c2",x"49",x"70",x"87"),
  2180 => (x"87",x"cf",x"05",x"99"),
  2181 => (x"bf",x"ec",x"d4",x"c2"),
  2182 => (x"6e",x"b9",x"ff",x"49"),
  2183 => (x"02",x"99",x"c1",x"99"),
  2184 => (x"cb",x"87",x"c0",x"c2"),
  2185 => (x"cf",x"cc",x"49",x"ee"),
  2186 => (x"58",x"a6",x"d0",x"87"),
  2187 => (x"d2",x"e8",x"49",x"c7"),
  2188 => (x"05",x"98",x"70",x"87"),
  2189 => (x"49",x"6e",x"87",x"c8"),
  2190 => (x"c1",x"02",x"99",x"c1"),
  2191 => (x"66",x"cc",x"87",x"c2"),
  2192 => (x"7e",x"bf",x"ec",x"4b"),
  2193 => (x"bf",x"f4",x"d4",x"c2"),
  2194 => (x"87",x"f5",x"e2",x"49"),
  2195 => (x"f3",x"cb",x"49",x"73"),
  2196 => (x"02",x"98",x"70",x"87"),
  2197 => (x"d4",x"c2",x"87",x"d7"),
  2198 => (x"c1",x"49",x"bf",x"d4"),
  2199 => (x"d8",x"d4",x"c2",x"b9"),
  2200 => (x"da",x"fd",x"71",x"59"),
  2201 => (x"49",x"ee",x"cb",x"87"),
  2202 => (x"70",x"87",x"cd",x"cb"),
  2203 => (x"e7",x"49",x"c7",x"4b"),
  2204 => (x"98",x"70",x"87",x"d1"),
  2205 => (x"87",x"c9",x"ff",x"05"),
  2206 => (x"99",x"c1",x"49",x"6e"),
  2207 => (x"87",x"c1",x"ff",x"05"),
  2208 => (x"bf",x"f4",x"d4",x"c2"),
  2209 => (x"c2",x"ba",x"c1",x"4a"),
  2210 => (x"fc",x"5a",x"f8",x"d4"),
  2211 => (x"c1",x"0a",x"7a",x"0a"),
  2212 => (x"a2",x"c0",x"c1",x"9a"),
  2213 => (x"87",x"fb",x"e8",x"49"),
  2214 => (x"e6",x"49",x"da",x"c1"),
  2215 => (x"a6",x"c8",x"87",x"e5"),
  2216 => (x"c2",x"78",x"c1",x"48"),
  2217 => (x"6e",x"48",x"ec",x"d4"),
  2218 => (x"f4",x"d4",x"c2",x"78"),
  2219 => (x"c7",x"c1",x"05",x"bf"),
  2220 => (x"c0",x"c0",x"c8",x"87"),
  2221 => (x"e0",x"d5",x"c2",x"4b"),
  2222 => (x"49",x"15",x"4d",x"7e"),
  2223 => (x"87",x"c3",x"e6",x"49"),
  2224 => (x"c0",x"02",x"98",x"70"),
  2225 => (x"b4",x"73",x"87",x"c2"),
  2226 => (x"05",x"2b",x"b7",x"c1"),
  2227 => (x"74",x"87",x"eb",x"ff"),
  2228 => (x"99",x"ff",x"c3",x"49"),
  2229 => (x"49",x"c0",x"1e",x"71"),
  2230 => (x"74",x"87",x"d5",x"fb"),
  2231 => (x"29",x"b7",x"c8",x"49"),
  2232 => (x"49",x"c1",x"1e",x"71"),
  2233 => (x"c8",x"87",x"c9",x"fb"),
  2234 => (x"49",x"fd",x"c3",x"86"),
  2235 => (x"c3",x"87",x"d4",x"e5"),
  2236 => (x"ce",x"e5",x"49",x"fa"),
  2237 => (x"87",x"d1",x"c8",x"87"),
  2238 => (x"ff",x"c3",x"49",x"74"),
  2239 => (x"2c",x"b7",x"c8",x"99"),
  2240 => (x"9c",x"74",x"b4",x"71"),
  2241 => (x"ff",x"87",x"df",x"02"),
  2242 => (x"49",x"7e",x"bf",x"c8"),
  2243 => (x"bf",x"f0",x"d4",x"c2"),
  2244 => (x"a9",x"e0",x"c2",x"89"),
  2245 => (x"87",x"c5",x"c0",x"03"),
  2246 => (x"cf",x"c0",x"4c",x"c0"),
  2247 => (x"f0",x"d4",x"c2",x"87"),
  2248 => (x"c0",x"78",x"6e",x"48"),
  2249 => (x"d4",x"c2",x"87",x"c6"),
  2250 => (x"78",x"c0",x"48",x"f0"),
  2251 => (x"99",x"c8",x"49",x"74"),
  2252 => (x"87",x"ce",x"c0",x"05"),
  2253 => (x"e4",x"49",x"f5",x"c3"),
  2254 => (x"49",x"70",x"87",x"c9"),
  2255 => (x"c0",x"02",x"99",x"c2"),
  2256 => (x"e8",x"c2",x"87",x"ea"),
  2257 => (x"c0",x"02",x"bf",x"ec"),
  2258 => (x"c1",x"48",x"87",x"ca"),
  2259 => (x"f0",x"e8",x"c2",x"88"),
  2260 => (x"87",x"d3",x"c0",x"58"),
  2261 => (x"c1",x"48",x"66",x"c4"),
  2262 => (x"7e",x"70",x"80",x"e0"),
  2263 => (x"c0",x"02",x"bf",x"6e"),
  2264 => (x"ff",x"4b",x"87",x"c5"),
  2265 => (x"c8",x"0f",x"73",x"49"),
  2266 => (x"78",x"c1",x"48",x"a6"),
  2267 => (x"99",x"c4",x"49",x"74"),
  2268 => (x"87",x"ce",x"c0",x"05"),
  2269 => (x"e3",x"49",x"f2",x"c3"),
  2270 => (x"49",x"70",x"87",x"c9"),
  2271 => (x"c0",x"02",x"99",x"c2"),
  2272 => (x"e8",x"c2",x"87",x"f0"),
  2273 => (x"48",x"7e",x"bf",x"ec"),
  2274 => (x"03",x"a8",x"b7",x"c7"),
  2275 => (x"6e",x"87",x"cb",x"c0"),
  2276 => (x"c2",x"80",x"c1",x"48"),
  2277 => (x"c0",x"58",x"f0",x"e8"),
  2278 => (x"66",x"c4",x"87",x"d3"),
  2279 => (x"80",x"e0",x"c1",x"48"),
  2280 => (x"bf",x"6e",x"7e",x"70"),
  2281 => (x"87",x"c5",x"c0",x"02"),
  2282 => (x"73",x"49",x"fe",x"4b"),
  2283 => (x"48",x"a6",x"c8",x"0f"),
  2284 => (x"fd",x"c3",x"78",x"c1"),
  2285 => (x"87",x"cb",x"e2",x"49"),
  2286 => (x"99",x"c2",x"49",x"70"),
  2287 => (x"87",x"e6",x"c0",x"02"),
  2288 => (x"bf",x"ec",x"e8",x"c2"),
  2289 => (x"87",x"c9",x"c0",x"02"),
  2290 => (x"48",x"ec",x"e8",x"c2"),
  2291 => (x"d0",x"c0",x"78",x"c0"),
  2292 => (x"4a",x"66",x"c4",x"87"),
  2293 => (x"6a",x"82",x"e0",x"c1"),
  2294 => (x"87",x"c5",x"c0",x"02"),
  2295 => (x"73",x"49",x"fd",x"4b"),
  2296 => (x"48",x"a6",x"c8",x"0f"),
  2297 => (x"fa",x"c3",x"78",x"c1"),
  2298 => (x"87",x"d7",x"e1",x"49"),
  2299 => (x"99",x"c2",x"49",x"70"),
  2300 => (x"87",x"ed",x"c0",x"02"),
  2301 => (x"bf",x"ec",x"e8",x"c2"),
  2302 => (x"a8",x"b7",x"c7",x"48"),
  2303 => (x"87",x"c9",x"c0",x"03"),
  2304 => (x"48",x"ec",x"e8",x"c2"),
  2305 => (x"d3",x"c0",x"78",x"c7"),
  2306 => (x"48",x"66",x"c4",x"87"),
  2307 => (x"70",x"80",x"e0",x"c1"),
  2308 => (x"02",x"bf",x"6e",x"7e"),
  2309 => (x"4b",x"87",x"c5",x"c0"),
  2310 => (x"0f",x"73",x"49",x"fc"),
  2311 => (x"c1",x"48",x"a6",x"c8"),
  2312 => (x"c3",x"48",x"74",x"78"),
  2313 => (x"7e",x"70",x"98",x"f0"),
  2314 => (x"c0",x"05",x"98",x"48"),
  2315 => (x"da",x"c1",x"87",x"ce"),
  2316 => (x"87",x"cf",x"e0",x"49"),
  2317 => (x"99",x"c2",x"49",x"70"),
  2318 => (x"87",x"d0",x"c2",x"02"),
  2319 => (x"c3",x"49",x"ee",x"cb"),
  2320 => (x"a6",x"d0",x"87",x"f6"),
  2321 => (x"e4",x"e8",x"c2",x"58"),
  2322 => (x"c2",x"50",x"c0",x"48"),
  2323 => (x"bf",x"97",x"e4",x"e8"),
  2324 => (x"87",x"d8",x"c1",x"05"),
  2325 => (x"cd",x"c0",x"05",x"6e"),
  2326 => (x"49",x"da",x"c1",x"87"),
  2327 => (x"87",x"e3",x"df",x"ff"),
  2328 => (x"c1",x"02",x"98",x"70"),
  2329 => (x"bf",x"e8",x"87",x"c6"),
  2330 => (x"ff",x"c3",x"49",x"4b"),
  2331 => (x"2b",x"b7",x"c8",x"99"),
  2332 => (x"d4",x"c2",x"b3",x"71"),
  2333 => (x"ff",x"49",x"bf",x"f4"),
  2334 => (x"cc",x"87",x"c6",x"da"),
  2335 => (x"c3",x"c3",x"49",x"66"),
  2336 => (x"02",x"98",x"70",x"87"),
  2337 => (x"c2",x"87",x"c6",x"c0"),
  2338 => (x"c1",x"48",x"e4",x"e8"),
  2339 => (x"e4",x"e8",x"c2",x"50"),
  2340 => (x"c0",x"05",x"bf",x"97"),
  2341 => (x"49",x"73",x"87",x"d6"),
  2342 => (x"05",x"99",x"f0",x"c3"),
  2343 => (x"c1",x"87",x"c7",x"ff"),
  2344 => (x"de",x"ff",x"49",x"da"),
  2345 => (x"98",x"70",x"87",x"dd"),
  2346 => (x"87",x"fa",x"fe",x"05"),
  2347 => (x"c2",x"48",x"a6",x"cc"),
  2348 => (x"78",x"bf",x"ec",x"e8"),
  2349 => (x"cc",x"49",x"66",x"cc"),
  2350 => (x"48",x"66",x"c4",x"91"),
  2351 => (x"7e",x"70",x"80",x"71"),
  2352 => (x"c0",x"02",x"bf",x"6e"),
  2353 => (x"cc",x"4b",x"87",x"c6"),
  2354 => (x"0f",x"73",x"49",x"66"),
  2355 => (x"c0",x"02",x"9d",x"75"),
  2356 => (x"02",x"6d",x"87",x"e9"),
  2357 => (x"6d",x"87",x"e4",x"c0"),
  2358 => (x"e6",x"dd",x"ff",x"49"),
  2359 => (x"c1",x"49",x"70",x"87"),
  2360 => (x"cb",x"c0",x"02",x"99"),
  2361 => (x"4b",x"a5",x"c4",x"87"),
  2362 => (x"bf",x"ec",x"e8",x"c2"),
  2363 => (x"0f",x"4b",x"6b",x"49"),
  2364 => (x"c0",x"02",x"85",x"c8"),
  2365 => (x"05",x"6d",x"87",x"c5"),
  2366 => (x"c8",x"87",x"dc",x"ff"),
  2367 => (x"c8",x"c0",x"02",x"66"),
  2368 => (x"ec",x"e8",x"c2",x"87"),
  2369 => (x"cf",x"f0",x"49",x"bf"),
  2370 => (x"26",x"8e",x"f0",x"87"),
  2371 => (x"26",x"4c",x"26",x"4d"),
  2372 => (x"00",x"4f",x"26",x"4b"),
  2373 => (x"00",x"00",x"00",x"00"),
  2374 => (x"00",x"00",x"00",x"10"),
  2375 => (x"14",x"11",x"12",x"58"),
  2376 => (x"23",x"1c",x"1b",x"1d"),
  2377 => (x"94",x"91",x"59",x"5a"),
  2378 => (x"f4",x"eb",x"f2",x"f5"),
  2379 => (x"00",x"00",x"00",x"00"),
  2380 => (x"00",x"00",x"00",x"00"),
  2381 => (x"00",x"00",x"00",x"00"),
  2382 => (x"ff",x"4a",x"71",x"1e"),
  2383 => (x"72",x"49",x"bf",x"c8"),
  2384 => (x"4f",x"26",x"48",x"a1"),
  2385 => (x"bf",x"c8",x"ff",x"1e"),
  2386 => (x"c0",x"c0",x"fe",x"89"),
  2387 => (x"a9",x"c0",x"c0",x"c0"),
  2388 => (x"c0",x"87",x"c4",x"01"),
  2389 => (x"c1",x"87",x"c2",x"4a"),
  2390 => (x"26",x"48",x"72",x"4a"),
  2391 => (x"00",x"00",x"00",x"4f"),
  2392 => (x"11",x"14",x"12",x"58"),
  2393 => (x"23",x"1c",x"1b",x"1d"),
  2394 => (x"91",x"94",x"59",x"5a"),
  2395 => (x"f4",x"eb",x"f2",x"f5"),
  2396 => (x"00",x"00",x"25",x"74"),
  2397 => (x"4f",x"54",x"55",x"41"),
  2398 => (x"54",x"4f",x"4f",x"42"),
  2399 => (x"17",x"00",x"42",x"47"),
  2400 => (x"17",x"00",x"00",x"1a"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

