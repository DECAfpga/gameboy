library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"f4e8c287",
    12 => x"48c0c84e",
    13 => x"d5c128c2",
    14 => x"ead6e5ea",
    15 => x"c1467149",
    16 => x"87f90188",
    17 => x"49f4e8c2",
    18 => x"48c4d6c2",
    19 => x"0389d089",
    20 => x"404040c0",
    21 => x"d087f640",
    22 => x"50c00581",
    23 => x"f90589c1",
    24 => x"c3d6c287",
    25 => x"ffd5c24d",
    26 => x"02ad744c",
    27 => x"0f2487c4",
    28 => x"e2c187f7",
    29 => x"d6c287d8",
    30 => x"d6c24dc3",
    31 => x"ad744cc3",
    32 => x"c487c602",
    33 => x"f50f6c8c",
    34 => x"87fd0087",
    35 => x"7186fc1e",
    36 => x"49c0ff4a",
    37 => x"c0c44869",
    38 => x"487e7098",
    39 => x"87f40298",
    40 => x"fc487972",
    41 => x"0e4f268e",
    42 => x"0e5c5b5e",
    43 => x"4cc04b71",
    44 => x"029a4a13",
    45 => x"497287cd",
    46 => x"c187d1ff",
    47 => x"9a4a1384",
    48 => x"7487f305",
    49 => x"264c2648",
    50 => x"1e4f264b",
    51 => x"1e731e72",
    52 => x"02114812",
    53 => x"c34b87ca",
    54 => x"739b98df",
    55 => x"87f00288",
    56 => x"4a264b26",
    57 => x"731e4f26",
    58 => x"c11e721e",
    59 => x"87ca048b",
    60 => x"02114812",
    61 => x"028887c4",
    62 => x"4a2687f1",
    63 => x"4f264b26",
    64 => x"731e741e",
    65 => x"c11e721e",
    66 => x"87cf048b",
    67 => x"02114812",
    68 => x"df4c87c9",
    69 => x"88749c98",
    70 => x"2687ec02",
    71 => x"264b264a",
    72 => x"1e4f264c",
    73 => x"73814873",
    74 => x"87c502a9",
    75 => x"f6055312",
    76 => x"0e4f2687",
    77 => x"0e5c5b5e",
    78 => x"d4ff4a71",
    79 => x"4b66cc4c",
    80 => x"718bc149",
    81 => x"87ce0299",
    82 => x"6c7cffc3",
    83 => x"c1497352",
    84 => x"0599718b",
    85 => x"4c2687f2",
    86 => x"4f264b26",
    87 => x"ff1e731e",
    88 => x"ffc34bd4",
    89 => x"c34a6b7b",
    90 => x"496b7bff",
    91 => x"b17232c8",
    92 => x"6b7bffc3",
    93 => x"7131c84a",
    94 => x"7bffc3b2",
    95 => x"32c8496b",
    96 => x"4871b172",
    97 => x"4f264b26",
    98 => x"5c5b5e0e",
    99 => x"4d710e5d",
   100 => x"754cd4ff",
   101 => x"98ffc348",
   102 => x"d6c27c70",
   103 => x"c805bfc4",
   104 => x"4866d087",
   105 => x"a6d430c9",
   106 => x"4966d058",
   107 => x"487129d8",
   108 => x"7098ffc3",
   109 => x"4966d07c",
   110 => x"487129d0",
   111 => x"7098ffc3",
   112 => x"4966d07c",
   113 => x"487129c8",
   114 => x"7098ffc3",
   115 => x"4866d07c",
   116 => x"7098ffc3",
   117 => x"d049757c",
   118 => x"c3487129",
   119 => x"7c7098ff",
   120 => x"f0c94b6c",
   121 => x"ffc34aff",
   122 => x"87cf05ab",
   123 => x"6c7c7149",
   124 => x"028ac14b",
   125 => x"ab7187c5",
   126 => x"7387f202",
   127 => x"264d2648",
   128 => x"264b264c",
   129 => x"49c01e4f",
   130 => x"c348d4ff",
   131 => x"81c178ff",
   132 => x"a9b7c8c3",
   133 => x"2687f104",
   134 => x"5b5e0e4f",
   135 => x"c00e5d5c",
   136 => x"f7c1f0ff",
   137 => x"c0c0c14d",
   138 => x"4bc0c0c0",
   139 => x"c487d6ff",
   140 => x"c04cdff8",
   141 => x"fd49751e",
   142 => x"86c487ce",
   143 => x"c005a8c1",
   144 => x"d4ff87e5",
   145 => x"78ffc348",
   146 => x"e1c01e73",
   147 => x"49e9c1f0",
   148 => x"c487f5fc",
   149 => x"05987086",
   150 => x"d4ff87ca",
   151 => x"78ffc348",
   152 => x"87cb48c1",
   153 => x"c187defe",
   154 => x"c6ff058c",
   155 => x"2648c087",
   156 => x"264c264d",
   157 => x"0e4f264b",
   158 => x"0e5c5b5e",
   159 => x"c1f0ffc0",
   160 => x"d4ff4cc1",
   161 => x"78ffc348",
   162 => x"f849fcca",
   163 => x"4bd387d9",
   164 => x"49741ec0",
   165 => x"c487f1fb",
   166 => x"05987086",
   167 => x"d4ff87ca",
   168 => x"78ffc348",
   169 => x"87cb48c1",
   170 => x"c187dafd",
   171 => x"dfff058b",
   172 => x"2648c087",
   173 => x"264b264c",
   174 => x"0000004f",
   175 => x"00444d43",
   176 => x"43484453",
   177 => x"69616620",
   178 => x"000a216c",
   179 => x"52524549",
   180 => x"00000000",
   181 => x"00495053",
   182 => x"74697257",
   183 => x"61662065",
   184 => x"64656c69",
   185 => x"5e0e000a",
   186 => x"0e5d5c5b",
   187 => x"ff4dffc3",
   188 => x"d0fc4bd4",
   189 => x"1eeac687",
   190 => x"c1f0e1c0",
   191 => x"c7fa49c8",
   192 => x"c186c487",
   193 => x"87c802a8",
   194 => x"c087ecfd",
   195 => x"87e8c148",
   196 => x"7087c9f9",
   197 => x"ffffcf49",
   198 => x"a9eac699",
   199 => x"fd87c802",
   200 => x"48c087d5",
   201 => x"7587d1c1",
   202 => x"4cf1c07b",
   203 => x"7087eafb",
   204 => x"ecc00298",
   205 => x"c01ec087",
   206 => x"fac1f0ff",
   207 => x"87c8f949",
   208 => x"987086c4",
   209 => x"7587da05",
   210 => x"75496b7b",
   211 => x"757b757b",
   212 => x"c17b757b",
   213 => x"c40299c0",
   214 => x"db48c187",
   215 => x"d748c087",
   216 => x"05acc287",
   217 => x"c0cb87ca",
   218 => x"87fbf449",
   219 => x"87c848c0",
   220 => x"fe058cc1",
   221 => x"48c087f6",
   222 => x"4c264d26",
   223 => x"4f264b26",
   224 => x"5c5b5e0e",
   225 => x"d0ff0e5d",
   226 => x"d0e5c04d",
   227 => x"c24cc0c1",
   228 => x"c148c4d6",
   229 => x"49d4cb78",
   230 => x"c787ccf4",
   231 => x"f97dc24b",
   232 => x"7dc387e3",
   233 => x"49741ec0",
   234 => x"c487ddf7",
   235 => x"05a8c186",
   236 => x"c24b87c1",
   237 => x"87cb05ab",
   238 => x"f349cccb",
   239 => x"48c087e9",
   240 => x"c187f6c0",
   241 => x"d4ff058b",
   242 => x"87dafc87",
   243 => x"58c8d6c2",
   244 => x"cd059870",
   245 => x"c01ec187",
   246 => x"d0c1f0ff",
   247 => x"87e8f649",
   248 => x"d4ff86c4",
   249 => x"78ffc348",
   250 => x"c287c3c3",
   251 => x"c258ccd6",
   252 => x"48d4ff7d",
   253 => x"c178ffc3",
   254 => x"264d2648",
   255 => x"264b264c",
   256 => x"5b5e0e4f",
   257 => x"fc0e5d5c",
   258 => x"ff4b7186",
   259 => x"7ec04cd4",
   260 => x"dfcdeec5",
   261 => x"7cffc34a",
   262 => x"fec3486c",
   263 => x"f8c005a8",
   264 => x"734d7487",
   265 => x"87cc029b",
   266 => x"731e66d4",
   267 => x"87c3f449",
   268 => x"87d486c4",
   269 => x"c448d0ff",
   270 => x"66d478d1",
   271 => x"7dffc34a",
   272 => x"f8058ac1",
   273 => x"5aa6d887",
   274 => x"7c7cffc3",
   275 => x"c5059b73",
   276 => x"48d0ff87",
   277 => x"4ac178d0",
   278 => x"058ac17e",
   279 => x"6e87f6fe",
   280 => x"268efc48",
   281 => x"264c264d",
   282 => x"1e4f264b",
   283 => x"4a711e73",
   284 => x"d4ff4bc0",
   285 => x"78ffc348",
   286 => x"c448d0ff",
   287 => x"d4ff78c3",
   288 => x"78ffc348",
   289 => x"ffc01e72",
   290 => x"49d1c1f0",
   291 => x"c487f9f3",
   292 => x"05987086",
   293 => x"c0c887d2",
   294 => x"4966cc1e",
   295 => x"c487e2fd",
   296 => x"ff4b7086",
   297 => x"78c248d0",
   298 => x"4b264873",
   299 => x"5e0e4f26",
   300 => x"0e5d5c5b",
   301 => x"ffc01ec0",
   302 => x"49c9c1f0",
   303 => x"d287c9f3",
   304 => x"d4d6c21e",
   305 => x"87f9fc49",
   306 => x"4cc086c8",
   307 => x"b7d284c1",
   308 => x"87f804ac",
   309 => x"97d4d6c2",
   310 => x"c0c349bf",
   311 => x"a9c0c199",
   312 => x"87e7c005",
   313 => x"97dbd6c2",
   314 => x"31d049bf",
   315 => x"97dcd6c2",
   316 => x"32c84abf",
   317 => x"d6c2b172",
   318 => x"4abf97dd",
   319 => x"cf4c71b1",
   320 => x"9cffffff",
   321 => x"34ca84c1",
   322 => x"c287e7c1",
   323 => x"bf97ddd6",
   324 => x"c631c149",
   325 => x"ded6c299",
   326 => x"c74abf97",
   327 => x"b1722ab7",
   328 => x"97d9d6c2",
   329 => x"cf4d4abf",
   330 => x"dad6c29d",
   331 => x"c34abf97",
   332 => x"c232ca9a",
   333 => x"bf97dbd6",
   334 => x"7333c24b",
   335 => x"dcd6c2b2",
   336 => x"c34bbf97",
   337 => x"b7c69bc0",
   338 => x"c2b2732b",
   339 => x"7148c181",
   340 => x"c1497030",
   341 => x"70307548",
   342 => x"c14c724d",
   343 => x"c8947184",
   344 => x"06adb7c0",
   345 => x"34c187cc",
   346 => x"c0c82db7",
   347 => x"ff01adb7",
   348 => x"487487f4",
   349 => x"4c264d26",
   350 => x"4f264b26",
   351 => x"5c5b5e0e",
   352 => x"86f80e5d",
   353 => x"48fcdec2",
   354 => x"d6c278c0",
   355 => x"49c01ef4",
   356 => x"c487d8fb",
   357 => x"05987086",
   358 => x"48c087c5",
   359 => x"c087f1c8",
   360 => x"c27ec14d",
   361 => x"df4aead7",
   362 => x"4bc849e8",
   363 => x"7087f7ec",
   364 => x"87c20598",
   365 => x"d8c27ec0",
   366 => x"f4df4ac6",
   367 => x"ec4bc849",
   368 => x"987087e4",
   369 => x"c087c205",
   370 => x"c0026e7e",
   371 => x"ddc287fd",
   372 => x"c24dbffa",
   373 => x"bf9ff2de",
   374 => x"d6c5487e",
   375 => x"c705a8ea",
   376 => x"faddc287",
   377 => x"87ce4dbf",
   378 => x"e9ca486e",
   379 => x"c502a8d5",
   380 => x"c748c087",
   381 => x"d6c287da",
   382 => x"49751ef4",
   383 => x"c487ecf9",
   384 => x"05987086",
   385 => x"48c087c5",
   386 => x"c287c5c7",
   387 => x"c04ac6d8",
   388 => x"c849c0e0",
   389 => x"87ceeb4b",
   390 => x"c8059870",
   391 => x"fcdec287",
   392 => x"d778c148",
   393 => x"ead7c287",
   394 => x"cce0c04a",
   395 => x"ea4bc849",
   396 => x"987087f4",
   397 => x"c087c502",
   398 => x"87d4c648",
   399 => x"97f2dec2",
   400 => x"d5c149bf",
   401 => x"87cd05a9",
   402 => x"97f3dec2",
   403 => x"eac249bf",
   404 => x"c5c002a9",
   405 => x"c548c087",
   406 => x"d6c287f6",
   407 => x"7ebf97f4",
   408 => x"a8e9c348",
   409 => x"87cec002",
   410 => x"ebc3486e",
   411 => x"c5c002a8",
   412 => x"c548c087",
   413 => x"d6c287da",
   414 => x"49bf97ff",
   415 => x"ccc00599",
   416 => x"c0d7c287",
   417 => x"c249bf97",
   418 => x"c5c002a9",
   419 => x"c448c087",
   420 => x"d7c287fe",
   421 => x"48bf97c1",
   422 => x"58f8dec2",
   423 => x"c1484c70",
   424 => x"fcdec288",
   425 => x"c2d7c258",
   426 => x"7549bf97",
   427 => x"c3d7c281",
   428 => x"c84abf97",
   429 => x"7ea17232",
   430 => x"48cce3c2",
   431 => x"d7c2786e",
   432 => x"48bf97c4",
   433 => x"c258a6c8",
   434 => x"02bffcde",
   435 => x"c287ccc2",
   436 => x"df4ac6d8",
   437 => x"4bc849dc",
   438 => x"7087cbe8",
   439 => x"c5c00298",
   440 => x"c348c087",
   441 => x"dec287ea",
   442 => x"c24cbff4",
   443 => x"c25ce0e3",
   444 => x"bf97d9d7",
   445 => x"c231c849",
   446 => x"bf97d8d7",
   447 => x"c249a14a",
   448 => x"bf97dad7",
   449 => x"7232d04a",
   450 => x"d7c249a1",
   451 => x"4abf97db",
   452 => x"a17232d8",
   453 => x"9166c449",
   454 => x"bfcce3c2",
   455 => x"d4e3c281",
   456 => x"e1d7c259",
   457 => x"c84abf97",
   458 => x"e0d7c232",
   459 => x"a24bbf97",
   460 => x"e2d7c24a",
   461 => x"d04bbf97",
   462 => x"4aa27333",
   463 => x"97e3d7c2",
   464 => x"9bcf4bbf",
   465 => x"a27333d8",
   466 => x"d8e3c24a",
   467 => x"748ac25a",
   468 => x"d8e3c292",
   469 => x"78a17248",
   470 => x"c287c1c1",
   471 => x"bf97c6d7",
   472 => x"c231c849",
   473 => x"bf97c5d7",
   474 => x"c549a14a",
   475 => x"81ffc731",
   476 => x"e3c229c9",
   477 => x"d7c259e0",
   478 => x"4abf97cb",
   479 => x"d7c232c8",
   480 => x"4bbf97ca",
   481 => x"66c44aa2",
   482 => x"c2826e92",
   483 => x"c25adce3",
   484 => x"c048d4e3",
   485 => x"d0e3c278",
   486 => x"78a17248",
   487 => x"48e0e3c2",
   488 => x"bfd4e3c2",
   489 => x"e4e3c278",
   490 => x"d8e3c248",
   491 => x"dec278bf",
   492 => x"c002bffc",
   493 => x"487487c9",
   494 => x"7e7030c4",
   495 => x"c287c9c0",
   496 => x"48bfdce3",
   497 => x"7e7030c4",
   498 => x"48c0dfc2",
   499 => x"48c1786e",
   500 => x"4d268ef8",
   501 => x"4b264c26",
   502 => x"00004f26",
   503 => x"33544146",
   504 => x"20202032",
   505 => x"00000000",
   506 => x"31544146",
   507 => x"20202036",
   508 => x"00000000",
   509 => x"33544146",
   510 => x"20202032",
   511 => x"00000000",
   512 => x"33544146",
   513 => x"20202032",
   514 => x"00000000",
   515 => x"31544146",
   516 => x"20202036",
   517 => x"00000000",
   518 => x"20202e2e",
   519 => x"20202020",
   520 => x"00202020",
   521 => x"5c5b5e0e",
   522 => x"4a710e5d",
   523 => x"bffcdec2",
   524 => x"7287cb02",
   525 => x"722bc74b",
   526 => x"9dffc14d",
   527 => x"4b7287c9",
   528 => x"4d722bc8",
   529 => x"c29dffc3",
   530 => x"83bfcce3",
   531 => x"bfc4f2c0",
   532 => x"87d902ab",
   533 => x"5bc8f2c0",
   534 => x"1ef4d6c2",
   535 => x"caf04973",
   536 => x"7086c487",
   537 => x"87c50598",
   538 => x"e6c048c0",
   539 => x"fcdec287",
   540 => x"87d202bf",
   541 => x"91c44975",
   542 => x"81f4d6c2",
   543 => x"ffcf4c69",
   544 => x"9cffffff",
   545 => x"497587cb",
   546 => x"d6c291c2",
   547 => x"699f81f4",
   548 => x"2648744c",
   549 => x"264c264d",
   550 => x"0e4f264b",
   551 => x"5d5c5b5e",
   552 => x"cc86f40e",
   553 => x"66c859a6",
   554 => x"7080c848",
   555 => x"78c0487e",
   556 => x"4949c11e",
   557 => x"c487d3c7",
   558 => x"9c4c7086",
   559 => x"87fac002",
   560 => x"4ac4dfc2",
   561 => x"e04966dc",
   562 => x"987087c1",
   563 => x"87eac002",
   564 => x"66dc4a74",
   565 => x"e04bcb49",
   566 => x"987087e6",
   567 => x"c087db02",
   568 => x"029c741e",
   569 => x"4dc087c4",
   570 => x"4dc187c2",
   571 => x"d9c64975",
   572 => x"7086c487",
   573 => x"ff059c4c",
   574 => x"9c7487c6",
   575 => x"87d7c102",
   576 => x"6e49a4dc",
   577 => x"da786948",
   578 => x"66c849a4",
   579 => x"c880c448",
   580 => x"699f58a6",
   581 => x"0866c448",
   582 => x"fcdec278",
   583 => x"87d202bf",
   584 => x"9f49a4d4",
   585 => x"ffc04969",
   586 => x"487199ff",
   587 => x"7e7030d0",
   588 => x"7ec087c2",
   589 => x"66c4486e",
   590 => x"66c480bf",
   591 => x"66c87808",
   592 => x"c878c048",
   593 => x"81cc4966",
   594 => x"79bf66c4",
   595 => x"d04966c8",
   596 => x"c179c081",
   597 => x"c087c248",
   598 => x"268ef448",
   599 => x"264c264d",
   600 => x"0e4f264b",
   601 => x"5d5c5b5e",
   602 => x"d04c710e",
   603 => x"6c4a4d66",
   604 => x"4da17249",
   605 => x"f8dec2b9",
   606 => x"baff4abf",
   607 => x"99719972",
   608 => x"87e4c002",
   609 => x"6b4ba4c4",
   610 => x"87d8fa49",
   611 => x"dec27b70",
   612 => x"6c49bff4",
   613 => x"757c7181",
   614 => x"f8dec2b9",
   615 => x"baff4abf",
   616 => x"99719972",
   617 => x"87dcff05",
   618 => x"4d267c75",
   619 => x"4b264c26",
   620 => x"731e4f26",
   621 => x"c24b711e",
   622 => x"49bfd0e3",
   623 => x"6a4aa3c4",
   624 => x"c28ac24a",
   625 => x"92bff4de",
   626 => x"c249a172",
   627 => x"4abff8de",
   628 => x"a1729a6b",
   629 => x"c8f2c049",
   630 => x"1e66c859",
   631 => x"87cbea71",
   632 => x"987086c4",
   633 => x"c087c405",
   634 => x"c187c248",
   635 => x"264b2648",
   636 => x"1e731e4f",
   637 => x"029b4b71",
   638 => x"c287e4c0",
   639 => x"735be4e3",
   640 => x"c28ac24a",
   641 => x"49bff4de",
   642 => x"d0e3c292",
   643 => x"807248bf",
   644 => x"58e8e3c2",
   645 => x"30c44871",
   646 => x"58c4dfc2",
   647 => x"c287edc0",
   648 => x"c248e0e3",
   649 => x"78bfd4e3",
   650 => x"48e4e3c2",
   651 => x"bfd8e3c2",
   652 => x"fcdec278",
   653 => x"87c902bf",
   654 => x"bff4dec2",
   655 => x"c731c449",
   656 => x"dce3c287",
   657 => x"31c449bf",
   658 => x"59c4dfc2",
   659 => x"4f264b26",
   660 => x"5c5b5e0e",
   661 => x"c04a710e",
   662 => x"029a724b",
   663 => x"da87e0c0",
   664 => x"699f49a2",
   665 => x"fcdec24b",
   666 => x"87cf02bf",
   667 => x"9f49a2d4",
   668 => x"c04c4969",
   669 => x"d09cffff",
   670 => x"c087c234",
   671 => x"73b3744c",
   672 => x"87edfd49",
   673 => x"4b264c26",
   674 => x"5e0e4f26",
   675 => x"0e5d5c5b",
   676 => x"a6c886f0",
   677 => x"ffffcf59",
   678 => x"c04cf8ff",
   679 => x"0266c47e",
   680 => x"d6c287d8",
   681 => x"78c048f0",
   682 => x"48e8d6c2",
   683 => x"bfe4e3c2",
   684 => x"ecd6c278",
   685 => x"e0e3c248",
   686 => x"dfc278bf",
   687 => x"50c048d1",
   688 => x"bfc0dfc2",
   689 => x"f0d6c249",
   690 => x"aa714abf",
   691 => x"87cbc403",
   692 => x"99cf4972",
   693 => x"87e9c005",
   694 => x"48c4f2c0",
   695 => x"bfe8d6c2",
   696 => x"f4d6c278",
   697 => x"e8d6c21e",
   698 => x"d6c249bf",
   699 => x"a1c148e8",
   700 => x"f6e57178",
   701 => x"c086c487",
   702 => x"c248c0f2",
   703 => x"cc78f4d6",
   704 => x"c0f2c087",
   705 => x"e0c048bf",
   706 => x"c4f2c080",
   707 => x"f0d6c258",
   708 => x"80c148bf",
   709 => x"58f4d6c2",
   710 => x"000c8027",
   711 => x"bf97bf00",
   712 => x"c2029d4d",
   713 => x"e5c387e5",
   714 => x"dec202ad",
   715 => x"c0f2c087",
   716 => x"a3cb4bbf",
   717 => x"cf4c1149",
   718 => x"d2c105ac",
   719 => x"df497587",
   720 => x"cd89c199",
   721 => x"c4dfc291",
   722 => x"4aa3c181",
   723 => x"a3c35112",
   724 => x"c551124a",
   725 => x"51124aa3",
   726 => x"124aa3c7",
   727 => x"4aa3c951",
   728 => x"a3ce5112",
   729 => x"d051124a",
   730 => x"51124aa3",
   731 => x"124aa3d2",
   732 => x"4aa3d451",
   733 => x"a3d65112",
   734 => x"d851124a",
   735 => x"51124aa3",
   736 => x"124aa3dc",
   737 => x"4aa3de51",
   738 => x"7ec15112",
   739 => x"7487fcc0",
   740 => x"0599c849",
   741 => x"7487edc0",
   742 => x"0599d049",
   743 => x"e0c087d3",
   744 => x"ccc00266",
   745 => x"c0497387",
   746 => x"700f66e0",
   747 => x"d3c00298",
   748 => x"c0056e87",
   749 => x"dfc287c6",
   750 => x"50c048c4",
   751 => x"bfc0f2c0",
   752 => x"87e9c248",
   753 => x"48d1dfc2",
   754 => x"c27e50c0",
   755 => x"49bfc0df",
   756 => x"bff0d6c2",
   757 => x"04aa714a",
   758 => x"cf87f5fb",
   759 => x"f8ffffff",
   760 => x"e4e3c24c",
   761 => x"c8c005bf",
   762 => x"fcdec287",
   763 => x"fac102bf",
   764 => x"ecd6c287",
   765 => x"ebf049bf",
   766 => x"f0d6c287",
   767 => x"48a6c458",
   768 => x"bfecd6c2",
   769 => x"fcdec278",
   770 => x"dbc002bf",
   771 => x"4966c487",
   772 => x"a9749974",
   773 => x"87c8c002",
   774 => x"c048a6c8",
   775 => x"87e7c078",
   776 => x"c148a6c8",
   777 => x"87dfc078",
   778 => x"cf4966c4",
   779 => x"a999f8ff",
   780 => x"87c8c002",
   781 => x"c048a6cc",
   782 => x"87c5c078",
   783 => x"c148a6cc",
   784 => x"48a6c878",
   785 => x"c87866cc",
   786 => x"dec00566",
   787 => x"4966c487",
   788 => x"dec289c2",
   789 => x"c291bff4",
   790 => x"48bfd0e3",
   791 => x"d6c28071",
   792 => x"d6c258ec",
   793 => x"78c048f0",
   794 => x"c087d5f9",
   795 => x"ffffcf48",
   796 => x"f04cf8ff",
   797 => x"264d268e",
   798 => x"264b264c",
   799 => x"0000004f",
   800 => x"00000000",
   801 => x"ffffffff",
   802 => x"48d4ff1e",
   803 => x"6878ffc3",
   804 => x"1e4f2648",
   805 => x"c348d4ff",
   806 => x"d0ff78ff",
   807 => x"78e1c048",
   808 => x"d448d4ff",
   809 => x"1e4f2678",
   810 => x"c048d0ff",
   811 => x"4f2678e0",
   812 => x"87d4ff1e",
   813 => x"02994970",
   814 => x"fbc087c6",
   815 => x"87f105a9",
   816 => x"4f264871",
   817 => x"5c5b5e0e",
   818 => x"c04b710e",
   819 => x"87f8fe4c",
   820 => x"02994970",
   821 => x"c087f9c0",
   822 => x"c002a9ec",
   823 => x"fbc087f2",
   824 => x"ebc002a9",
   825 => x"b766cc87",
   826 => x"87c703ac",
   827 => x"c20266d0",
   828 => x"71537187",
   829 => x"87c20299",
   830 => x"cbfe84c1",
   831 => x"99497087",
   832 => x"c087cd02",
   833 => x"c702a9ec",
   834 => x"a9fbc087",
   835 => x"87d5ff05",
   836 => x"c30266d0",
   837 => x"7b97c087",
   838 => x"05a9ecc0",
   839 => x"4a7487c4",
   840 => x"4a7487c5",
   841 => x"728a0ac0",
   842 => x"264c2648",
   843 => x"1e4f264b",
   844 => x"7087d5fd",
   845 => x"f0c04a49",
   846 => x"87c904aa",
   847 => x"01aaf9c0",
   848 => x"f0c087c3",
   849 => x"aac1c18a",
   850 => x"c187c904",
   851 => x"c301aada",
   852 => x"8af7c087",
   853 => x"4f264872",
   854 => x"5c5b5e0e",
   855 => x"86f80e5d",
   856 => x"7ec04c71",
   857 => x"c087ecfc",
   858 => x"f8f7c04b",
   859 => x"c049bf97",
   860 => x"87cf04a9",
   861 => x"c187f9fc",
   862 => x"f8f7c083",
   863 => x"ab49bf97",
   864 => x"c087f106",
   865 => x"bf97f8f7",
   866 => x"fb87cf02",
   867 => x"497087fa",
   868 => x"87c60299",
   869 => x"05a9ecc0",
   870 => x"4bc087f1",
   871 => x"7087e9fb",
   872 => x"87e4fb4d",
   873 => x"fb58a6c8",
   874 => x"4a7087de",
   875 => x"a4c883c1",
   876 => x"49699749",
   877 => x"87da05ad",
   878 => x"9749a4c9",
   879 => x"66c44969",
   880 => x"87ce05a9",
   881 => x"9749a4ca",
   882 => x"05aa4969",
   883 => x"7ec187c4",
   884 => x"ecc087d0",
   885 => x"87c602ad",
   886 => x"05adfbc0",
   887 => x"4bc087c4",
   888 => x"026e7ec1",
   889 => x"fa87f5fe",
   890 => x"487387fd",
   891 => x"4d268ef8",
   892 => x"4b264c26",
   893 => x"00004f26",
   894 => x"1e731e00",
   895 => x"c84bd4ff",
   896 => x"d0ff4a66",
   897 => x"78c5c848",
   898 => x"c148d4ff",
   899 => x"7b1178d4",
   900 => x"f9058ac1",
   901 => x"48d0ff87",
   902 => x"4b2678c4",
   903 => x"5e0e4f26",
   904 => x"0e5d5c5b",
   905 => x"7e7186f8",
   906 => x"e3c21e6e",
   907 => x"eae949f4",
   908 => x"7086c487",
   909 => x"e4c40298",
   910 => x"cce6c187",
   911 => x"496e4cbf",
   912 => x"c887d5fc",
   913 => x"987058a6",
   914 => x"c487c505",
   915 => x"78c148a6",
   916 => x"c548d0ff",
   917 => x"48d4ff78",
   918 => x"c478d5c1",
   919 => x"89c14966",
   920 => x"e6c131c6",
   921 => x"4abf97c4",
   922 => x"ffb07148",
   923 => x"ff7808d4",
   924 => x"78c448d0",
   925 => x"97f0e3c2",
   926 => x"99d049bf",
   927 => x"c587dd02",
   928 => x"48d4ff78",
   929 => x"c078d6c1",
   930 => x"48d4ff4a",
   931 => x"c178ffc3",
   932 => x"aae0c082",
   933 => x"ff87f204",
   934 => x"78c448d0",
   935 => x"c348d4ff",
   936 => x"d0ff78ff",
   937 => x"ff78c548",
   938 => x"d3c148d4",
   939 => x"ff78c178",
   940 => x"78c448d0",
   941 => x"06acb7c0",
   942 => x"c287cbc2",
   943 => x"4bbffce3",
   944 => x"737e748c",
   945 => x"ddc1029b",
   946 => x"4dc0c887",
   947 => x"abb7c08b",
   948 => x"c887c603",
   949 => x"c04da3c0",
   950 => x"f0e3c24b",
   951 => x"d049bf97",
   952 => x"87cf0299",
   953 => x"e3c21ec0",
   954 => x"c5eb49f4",
   955 => x"7086c487",
   956 => x"c287d84c",
   957 => x"c21ef4d6",
   958 => x"ea49f4e3",
   959 => x"4c7087f4",
   960 => x"d6c21e75",
   961 => x"f0fb49f4",
   962 => x"7486c887",
   963 => x"87c5059c",
   964 => x"cac148c0",
   965 => x"c21ec187",
   966 => x"e949f4e3",
   967 => x"86c487c5",
   968 => x"fe059b73",
   969 => x"4c6e87e3",
   970 => x"06acb7c0",
   971 => x"e3c287d1",
   972 => x"78c048f4",
   973 => x"78c080d0",
   974 => x"e4c280f4",
   975 => x"c078bfc0",
   976 => x"fd01acb7",
   977 => x"d0ff87f5",
   978 => x"ff78c548",
   979 => x"d3c148d4",
   980 => x"ff78c078",
   981 => x"78c448d0",
   982 => x"c2c048c1",
   983 => x"f848c087",
   984 => x"264d268e",
   985 => x"264b264c",
   986 => x"5b5e0e4f",
   987 => x"fc0e5d5c",
   988 => x"c04d7186",
   989 => x"04ad4c4b",
   990 => x"c087e8c0",
   991 => x"741ed8f5",
   992 => x"87c4029c",
   993 => x"87c24ac0",
   994 => x"49724ac1",
   995 => x"c487fbeb",
   996 => x"c17e7086",
   997 => x"c2056e83",
   998 => x"c14b7587",
   999 => x"06ab7584",
  1000 => x"6e87d8ff",
  1001 => x"268efc48",
  1002 => x"264c264d",
  1003 => x"1e4f264b",
  1004 => x"66c44a71",
  1005 => x"7287c505",
  1006 => x"87e2f949",
  1007 => x"5e0e4f26",
  1008 => x"0e5d5c5b",
  1009 => x"4c7186fc",
  1010 => x"c291de49",
  1011 => x"714de0e4",
  1012 => x"026d9785",
  1013 => x"c287dcc1",
  1014 => x"49bfd0e4",
  1015 => x"fe718174",
  1016 => x"7e7087c7",
  1017 => x"c0029848",
  1018 => x"e4c287f2",
  1019 => x"4a704bd4",
  1020 => x"c4ff49cb",
  1021 => x"4b7487ed",
  1022 => x"e6c193cc",
  1023 => x"83c483d0",
  1024 => x"7bc0c1c1",
  1025 => x"c4c14974",
  1026 => x"7b7587ce",
  1027 => x"97c8e6c1",
  1028 => x"c21e49bf",
  1029 => x"fe49d4e4",
  1030 => x"86c487d5",
  1031 => x"c3c14974",
  1032 => x"49c087f6",
  1033 => x"87d1c5c1",
  1034 => x"48ece3c2",
  1035 => x"c04950c0",
  1036 => x"fc87e6e2",
  1037 => x"264d268e",
  1038 => x"264b264c",
  1039 => x"0000004f",
  1040 => x"64616f4c",
  1041 => x"2e676e69",
  1042 => x"00002e2e",
  1043 => x"61422080",
  1044 => x"00006b63",
  1045 => x"64616f4c",
  1046 => x"202e2a20",
  1047 => x"00000000",
  1048 => x"0000203a",
  1049 => x"61422080",
  1050 => x"00006b63",
  1051 => x"78452080",
  1052 => x"00007469",
  1053 => x"49204453",
  1054 => x"2e74696e",
  1055 => x"0000002e",
  1056 => x"00004b4f",
  1057 => x"544f4f42",
  1058 => x"20202020",
  1059 => x"004d4f52",
  1060 => x"711e731e",
  1061 => x"e4c2494b",
  1062 => x"7181bfd0",
  1063 => x"7087cafb",
  1064 => x"c4029a4a",
  1065 => x"e7e64987",
  1066 => x"d0e4c287",
  1067 => x"7378c048",
  1068 => x"87fac149",
  1069 => x"4f264b26",
  1070 => x"711e731e",
  1071 => x"4aa3c44b",
  1072 => x"87d0c102",
  1073 => x"dc028ac1",
  1074 => x"c0028a87",
  1075 => x"058a87f2",
  1076 => x"c287d3c1",
  1077 => x"02bfd0e4",
  1078 => x"4887cbc1",
  1079 => x"e4c288c1",
  1080 => x"c1c158d4",
  1081 => x"d0e4c287",
  1082 => x"89c649bf",
  1083 => x"59d4e4c2",
  1084 => x"03a9b7c0",
  1085 => x"c287efc0",
  1086 => x"c048d0e4",
  1087 => x"87e6c078",
  1088 => x"bfcce4c2",
  1089 => x"c287df02",
  1090 => x"48bfd0e4",
  1091 => x"e4c280c1",
  1092 => x"87d258d4",
  1093 => x"bfcce4c2",
  1094 => x"c287cb02",
  1095 => x"48bfd0e4",
  1096 => x"e4c280c6",
  1097 => x"497358d4",
  1098 => x"4b2687c4",
  1099 => x"5e0e4f26",
  1100 => x"0e5d5c5b",
  1101 => x"a6d086f0",
  1102 => x"f4d6c259",
  1103 => x"c24cc04d",
  1104 => x"c148cce4",
  1105 => x"48a6c878",
  1106 => x"7e7578c0",
  1107 => x"bfd0e4c2",
  1108 => x"06a8c048",
  1109 => x"c887c0c1",
  1110 => x"7e755ca6",
  1111 => x"48f4d6c2",
  1112 => x"f2c00298",
  1113 => x"4d66c487",
  1114 => x"1ed8f5c0",
  1115 => x"c40266cc",
  1116 => x"c24cc087",
  1117 => x"744cc187",
  1118 => x"87cee449",
  1119 => x"7e7086c4",
  1120 => x"66c885c1",
  1121 => x"cc80c148",
  1122 => x"e4c258a6",
  1123 => x"03adbfd0",
  1124 => x"056e87c5",
  1125 => x"6e87d1ff",
  1126 => x"754cc04d",
  1127 => x"dcc3029d",
  1128 => x"d8f5c087",
  1129 => x"0266cc1e",
  1130 => x"a6c887c7",
  1131 => x"c578c048",
  1132 => x"48a6c887",
  1133 => x"66c878c1",
  1134 => x"87cee349",
  1135 => x"7e7086c4",
  1136 => x"c2029848",
  1137 => x"cb4987e4",
  1138 => x"49699781",
  1139 => x"c10299d0",
  1140 => x"497487d4",
  1141 => x"e6c191cc",
  1142 => x"c2c181d0",
  1143 => x"81c879d0",
  1144 => x"7451ffc3",
  1145 => x"c291de49",
  1146 => x"714de0e4",
  1147 => x"97c1c285",
  1148 => x"49a5c17d",
  1149 => x"c251e0c0",
  1150 => x"bf97c4df",
  1151 => x"c187d202",
  1152 => x"4ba5c284",
  1153 => x"4ac4dfc2",
  1154 => x"fcfe49db",
  1155 => x"d9c187d5",
  1156 => x"49a5cd87",
  1157 => x"84c151c0",
  1158 => x"6e4ba5c2",
  1159 => x"fe49cb4a",
  1160 => x"c187c0fc",
  1161 => x"497487c4",
  1162 => x"e6c191cc",
  1163 => x"fec081d0",
  1164 => x"dfc279fe",
  1165 => x"02bf97c4",
  1166 => x"497487d8",
  1167 => x"84c191de",
  1168 => x"4be0e4c2",
  1169 => x"dfc28371",
  1170 => x"49dd4ac4",
  1171 => x"87d3fbfe",
  1172 => x"4b7487d8",
  1173 => x"e4c293de",
  1174 => x"a3cb83e0",
  1175 => x"c151c049",
  1176 => x"4a6e7384",
  1177 => x"fafe49cb",
  1178 => x"66c887f9",
  1179 => x"cc80c148",
  1180 => x"acc758a6",
  1181 => x"87c5c003",
  1182 => x"e4fc056e",
  1183 => x"03acc787",
  1184 => x"c287e4c0",
  1185 => x"c048cce4",
  1186 => x"cc497478",
  1187 => x"d0e6c191",
  1188 => x"fefec081",
  1189 => x"de497479",
  1190 => x"e0e4c291",
  1191 => x"c151c081",
  1192 => x"04acc784",
  1193 => x"c187dcff",
  1194 => x"c048ece7",
  1195 => x"c180f750",
  1196 => x"c140d4cc",
  1197 => x"c878ccc1",
  1198 => x"f8c2c180",
  1199 => x"4966cc78",
  1200 => x"87d4f9c0",
  1201 => x"4d268ef0",
  1202 => x"4b264c26",
  1203 => x"731e4f26",
  1204 => x"494b711e",
  1205 => x"e6c191cc",
  1206 => x"a1c881d0",
  1207 => x"c4e6c14a",
  1208 => x"c9501248",
  1209 => x"f7c04aa1",
  1210 => x"501248f8",
  1211 => x"e6c181ca",
  1212 => x"501148c8",
  1213 => x"97c8e6c1",
  1214 => x"c01e49bf",
  1215 => x"87eff249",
  1216 => x"e9f84973",
  1217 => x"268efc87",
  1218 => x"1e4f264b",
  1219 => x"f9c049c0",
  1220 => x"4f2687e7",
  1221 => x"494a711e",
  1222 => x"e6c191cc",
  1223 => x"81c881d0",
  1224 => x"48ece3c2",
  1225 => x"f0c05011",
  1226 => x"f5fe49a2",
  1227 => x"49c087de",
  1228 => x"2687e6d6",
  1229 => x"d4ff1e4f",
  1230 => x"7affc34a",
  1231 => x"c048d0ff",
  1232 => x"7ade78e1",
  1233 => x"c8487a71",
  1234 => x"7a7028b7",
  1235 => x"b7d04871",
  1236 => x"717a7028",
  1237 => x"28b7d848",
  1238 => x"d0ff7a70",
  1239 => x"78e0c048",
  1240 => x"5e0e4f26",
  1241 => x"0e5d5c5b",
  1242 => x"4d7186f4",
  1243 => x"c191cc49",
  1244 => x"c881d0e6",
  1245 => x"a1ca4aa1",
  1246 => x"48a6c47e",
  1247 => x"bfe8e3c2",
  1248 => x"bf976e78",
  1249 => x"4c66c44b",
  1250 => x"48122c73",
  1251 => x"7058a6cc",
  1252 => x"c984c19c",
  1253 => x"49699781",
  1254 => x"c204acb7",
  1255 => x"6e4cc087",
  1256 => x"c84abf97",
  1257 => x"31724966",
  1258 => x"66c4b9ff",
  1259 => x"72487499",
  1260 => x"b14a7030",
  1261 => x"59ece3c2",
  1262 => x"87f9fd71",
  1263 => x"e4c21ec7",
  1264 => x"c11ebfc8",
  1265 => x"c21ed0e6",
  1266 => x"bf97ece3",
  1267 => x"87f4c149",
  1268 => x"f5c04975",
  1269 => x"8ee887c2",
  1270 => x"4c264d26",
  1271 => x"4f264b26",
  1272 => x"711e731e",
  1273 => x"f9fd494b",
  1274 => x"fd497387",
  1275 => x"4b2687f4",
  1276 => x"731e4f26",
  1277 => x"c24b711e",
  1278 => x"d6024aa3",
  1279 => x"058ac187",
  1280 => x"c287e2c0",
  1281 => x"02bfc8e4",
  1282 => x"c14887db",
  1283 => x"cce4c288",
  1284 => x"c287d258",
  1285 => x"02bfcce4",
  1286 => x"e4c287cb",
  1287 => x"c148bfc8",
  1288 => x"cce4c280",
  1289 => x"c21ec758",
  1290 => x"1ebfc8e4",
  1291 => x"1ed0e6c1",
  1292 => x"97ece3c2",
  1293 => x"87cc49bf",
  1294 => x"f3c04973",
  1295 => x"8ef487da",
  1296 => x"4f264b26",
  1297 => x"5c5b5e0e",
  1298 => x"ccff0e5d",
  1299 => x"a6e4c086",
  1300 => x"48a6cc59",
  1301 => x"80c478c0",
  1302 => x"80c478c0",
  1303 => x"7866c8c1",
  1304 => x"78c180c4",
  1305 => x"78c180c4",
  1306 => x"48cce4c2",
  1307 => x"e2e078c1",
  1308 => x"87fce087",
  1309 => x"7087d1e0",
  1310 => x"acfbc04c",
  1311 => x"87f3c102",
  1312 => x"0566e0c0",
  1313 => x"c187e8c1",
  1314 => x"c44a66c4",
  1315 => x"c17e6a82",
  1316 => x"6e48d4c1",
  1317 => x"20412049",
  1318 => x"c1511041",
  1319 => x"c14866c4",
  1320 => x"6a78cecb",
  1321 => x"7481c749",
  1322 => x"66c4c151",
  1323 => x"c181c849",
  1324 => x"48a6d851",
  1325 => x"c4c178c2",
  1326 => x"81c94966",
  1327 => x"c4c151c0",
  1328 => x"81ca4966",
  1329 => x"1ec151c0",
  1330 => x"496a1ed8",
  1331 => x"dfff81c8",
  1332 => x"86c887f2",
  1333 => x"4866c8c1",
  1334 => x"c701a8c0",
  1335 => x"48a6d087",
  1336 => x"87cf78c1",
  1337 => x"4866c8c1",
  1338 => x"a6d888c1",
  1339 => x"ff87c458",
  1340 => x"7487fdde",
  1341 => x"dacd029c",
  1342 => x"4866d087",
  1343 => x"a866ccc1",
  1344 => x"87cfcd03",
  1345 => x"c048a6c8",
  1346 => x"ddff7e78",
  1347 => x"4c7087fa",
  1348 => x"05acd0c1",
  1349 => x"c487e7c2",
  1350 => x"786e48a6",
  1351 => x"7087d0e0",
  1352 => x"66cc487e",
  1353 => x"87c506a8",
  1354 => x"6e48a6cc",
  1355 => x"d7ddff78",
  1356 => x"c04c7087",
  1357 => x"c105acec",
  1358 => x"66d087ee",
  1359 => x"c191cc49",
  1360 => x"c48166c4",
  1361 => x"4d6a4aa1",
  1362 => x"6e4aa1c8",
  1363 => x"d4ccc152",
  1364 => x"f3dcff79",
  1365 => x"9c4c7087",
  1366 => x"c087d902",
  1367 => x"d302acfb",
  1368 => x"ff557487",
  1369 => x"7087e1dc",
  1370 => x"c7029c4c",
  1371 => x"acfbc087",
  1372 => x"87edff05",
  1373 => x"c255e0c0",
  1374 => x"97c055c1",
  1375 => x"66e0c07d",
  1376 => x"a866c448",
  1377 => x"d087db05",
  1378 => x"66d44866",
  1379 => x"87ca04a8",
  1380 => x"c14866d0",
  1381 => x"58a6d480",
  1382 => x"66d487c8",
  1383 => x"d888c148",
  1384 => x"dbff58a6",
  1385 => x"4c7087e2",
  1386 => x"05acd0c1",
  1387 => x"66dc87c9",
  1388 => x"c080c148",
  1389 => x"c158a6e0",
  1390 => x"fd02acd0",
  1391 => x"486e87d9",
  1392 => x"a866e0c0",
  1393 => x"87ebc905",
  1394 => x"48a6e4c0",
  1395 => x"487478c0",
  1396 => x"c888fbc0",
  1397 => x"987058a6",
  1398 => x"87ddc902",
  1399 => x"c888cb48",
  1400 => x"987058a6",
  1401 => x"87cfc102",
  1402 => x"c888c948",
  1403 => x"987058a6",
  1404 => x"87ffc302",
  1405 => x"c888c448",
  1406 => x"987058a6",
  1407 => x"4887cf02",
  1408 => x"a6c888c1",
  1409 => x"02987058",
  1410 => x"c887e8c3",
  1411 => x"a6c887dc",
  1412 => x"78f0c048",
  1413 => x"87f0d9ff",
  1414 => x"ecc04c70",
  1415 => x"c3c002ac",
  1416 => x"5ca6cc87",
  1417 => x"02acecc0",
  1418 => x"d9ff87cd",
  1419 => x"4c7087da",
  1420 => x"05acecc0",
  1421 => x"c087f3ff",
  1422 => x"c002acec",
  1423 => x"d9ff87c4",
  1424 => x"1ec087c6",
  1425 => x"66d81eca",
  1426 => x"c191cc49",
  1427 => x"714866cc",
  1428 => x"58a6cc80",
  1429 => x"c44866c8",
  1430 => x"58a6d080",
  1431 => x"49bf66cc",
  1432 => x"87e0d9ff",
  1433 => x"1ede1ec1",
  1434 => x"49bf66d4",
  1435 => x"87d4d9ff",
  1436 => x"497086d0",
  1437 => x"8808c048",
  1438 => x"58a6ecc0",
  1439 => x"c006a8c0",
  1440 => x"e8c087ee",
  1441 => x"a8dd4866",
  1442 => x"87e4c003",
  1443 => x"49bf66c4",
  1444 => x"8166e8c0",
  1445 => x"c051e0c0",
  1446 => x"c14966e8",
  1447 => x"bf66c481",
  1448 => x"51c1c281",
  1449 => x"4966e8c0",
  1450 => x"66c481c2",
  1451 => x"51c081bf",
  1452 => x"cbc1486e",
  1453 => x"496e78ce",
  1454 => x"66d881c8",
  1455 => x"c9496e51",
  1456 => x"5166dc81",
  1457 => x"81ca496e",
  1458 => x"d85166c8",
  1459 => x"80c14866",
  1460 => x"d058a6dc",
  1461 => x"66d44866",
  1462 => x"cbc004a8",
  1463 => x"4866d087",
  1464 => x"a6d480c1",
  1465 => x"87d1c558",
  1466 => x"c14866d4",
  1467 => x"58a6d888",
  1468 => x"ff87c6c5",
  1469 => x"c087f8d8",
  1470 => x"ff58a6ec",
  1471 => x"c087f0d8",
  1472 => x"c058a6f0",
  1473 => x"c005a8ec",
  1474 => x"48a687c9",
  1475 => x"7866e8c0",
  1476 => x"ff87c4c0",
  1477 => x"d087f1d5",
  1478 => x"91cc4966",
  1479 => x"4866c4c1",
  1480 => x"a6c88071",
  1481 => x"4a66c458",
  1482 => x"66c482c8",
  1483 => x"c081ca49",
  1484 => x"c05166e8",
  1485 => x"c14966ec",
  1486 => x"66e8c081",
  1487 => x"7148c189",
  1488 => x"c1497030",
  1489 => x"7a977189",
  1490 => x"bfe8e3c2",
  1491 => x"66e8c049",
  1492 => x"4a6a9729",
  1493 => x"c0987148",
  1494 => x"c458a6f4",
  1495 => x"80c44866",
  1496 => x"c858a6cc",
  1497 => x"c04dbf66",
  1498 => x"6e4866e0",
  1499 => x"c5c002a8",
  1500 => x"c07ec087",
  1501 => x"7ec187c2",
  1502 => x"e0c01e6e",
  1503 => x"ff49751e",
  1504 => x"c887c1d5",
  1505 => x"c04c7086",
  1506 => x"c106acb7",
  1507 => x"857487d4",
  1508 => x"49bf66c8",
  1509 => x"7581e0c0",
  1510 => x"c1c14b89",
  1511 => x"fe714ae0",
  1512 => x"c287c0e6",
  1513 => x"c07e7585",
  1514 => x"c14866e4",
  1515 => x"a6e8c080",
  1516 => x"66f0c058",
  1517 => x"7081c149",
  1518 => x"c5c002a9",
  1519 => x"c04dc087",
  1520 => x"4dc187c2",
  1521 => x"66cc1e75",
  1522 => x"e0c049bf",
  1523 => x"8966c481",
  1524 => x"66c81e71",
  1525 => x"ebd3ff49",
  1526 => x"c086c887",
  1527 => x"ff01a8b7",
  1528 => x"e4c087c5",
  1529 => x"d3c00266",
  1530 => x"4966c487",
  1531 => x"e4c081c9",
  1532 => x"66c45166",
  1533 => x"e2cdc148",
  1534 => x"87cec078",
  1535 => x"c94966c4",
  1536 => x"c451c281",
  1537 => x"cfc14866",
  1538 => x"66d078e0",
  1539 => x"a866d448",
  1540 => x"87cbc004",
  1541 => x"c14866d0",
  1542 => x"58a6d480",
  1543 => x"d487dac0",
  1544 => x"88c14866",
  1545 => x"c058a6d8",
  1546 => x"d2ff87cf",
  1547 => x"4c7087c2",
  1548 => x"ff87c6c0",
  1549 => x"7087f9d1",
  1550 => x"4866dc4c",
  1551 => x"e0c080c1",
  1552 => x"9c7458a6",
  1553 => x"87cbc002",
  1554 => x"c14866d0",
  1555 => x"04a866cc",
  1556 => x"d087f1f2",
  1557 => x"a8c74866",
  1558 => x"87e1c003",
  1559 => x"c24c66d0",
  1560 => x"c048cce4",
  1561 => x"cc497478",
  1562 => x"66c4c191",
  1563 => x"4aa1c481",
  1564 => x"52c04a6a",
  1565 => x"c784c179",
  1566 => x"e2ff04ac",
  1567 => x"66e0c087",
  1568 => x"87e2c002",
  1569 => x"4966c4c1",
  1570 => x"c181d4c1",
  1571 => x"c14a66c4",
  1572 => x"52c082dc",
  1573 => x"79d4ccc1",
  1574 => x"4966c4c1",
  1575 => x"c181d8c1",
  1576 => x"c079e4c1",
  1577 => x"c4c187d6",
  1578 => x"d4c14966",
  1579 => x"66c4c181",
  1580 => x"82d8c14a",
  1581 => x"7aecc1c1",
  1582 => x"79cbccc1",
  1583 => x"4966c4c1",
  1584 => x"c181e0c1",
  1585 => x"ff79f2cf",
  1586 => x"cc87dccf",
  1587 => x"ccff4866",
  1588 => x"264d268e",
  1589 => x"264b264c",
  1590 => x"1ec71e4f",
  1591 => x"bfc8e4c2",
  1592 => x"d0e6c11e",
  1593 => x"ece3c21e",
  1594 => x"ed49bf97",
  1595 => x"e6c187d6",
  1596 => x"e1c049d0",
  1597 => x"8ef487f0",
  1598 => x"c11e4f26",
  1599 => x"c048c4e6",
  1600 => x"f0d5c250",
  1601 => x"d4ff49bf",
  1602 => x"48c087d4",
  1603 => x"731e4f26",
  1604 => x"87d9c71e",
  1605 => x"48d4e4c2",
  1606 => x"d4ff50c0",
  1607 => x"78ffc348",
  1608 => x"49f4c1c1",
  1609 => x"87ffddfe",
  1610 => x"87d4e9fe",
  1611 => x"cd029870",
  1612 => x"c7f1fe87",
  1613 => x"02987087",
  1614 => x"4ac187c4",
  1615 => x"4ac087c2",
  1616 => x"c8029a72",
  1617 => x"c0c2c187",
  1618 => x"daddfe49",
  1619 => x"c8e4c287",
  1620 => x"c278c048",
  1621 => x"c048ece3",
  1622 => x"fcfd4950",
  1623 => x"87dafe87",
  1624 => x"029b4b70",
  1625 => x"e7c187cf",
  1626 => x"49c75bec",
  1627 => x"c187e9de",
  1628 => x"c4e0c049",
  1629 => x"87efc287",
  1630 => x"87e5e1c0",
  1631 => x"4b2687fa",
  1632 => x"00004f26",
  1633 => x"00000000",
  1634 => x"00000000",
  1635 => x"00000001",
  1636 => x"00000fbe",
  1637 => x"00002920",
  1638 => x"00000000",
  1639 => x"00000fbe",
  1640 => x"0000293e",
  1641 => x"00000000",
  1642 => x"00000fbe",
  1643 => x"0000295c",
  1644 => x"00000000",
  1645 => x"00000fbe",
  1646 => x"0000297a",
  1647 => x"00000000",
  1648 => x"00000fbe",
  1649 => x"00002998",
  1650 => x"00000000",
  1651 => x"00000fbe",
  1652 => x"000029b6",
  1653 => x"00000000",
  1654 => x"00000fbe",
  1655 => x"000029d4",
  1656 => x"00000000",
  1657 => x"00001314",
  1658 => x"00000000",
  1659 => x"00000000",
  1660 => x"000010b8",
  1661 => x"00000000",
  1662 => x"00000000",
  1663 => x"00001084",
  1664 => x"db86fc1e",
  1665 => x"fc7e7087",
  1666 => x"1e4f268e",
  1667 => x"c048f0fe",
  1668 => x"7909cd78",
  1669 => x"1e4f2609",
  1670 => x"49c0e8c1",
  1671 => x"4f2687ed",
  1672 => x"bff0fe1e",
  1673 => x"1e4f2648",
  1674 => x"c148f0fe",
  1675 => x"1e4f2678",
  1676 => x"c048f0fe",
  1677 => x"1e4f2678",
  1678 => x"52c04a71",
  1679 => x"0e4f2651",
  1680 => x"5d5c5b5e",
  1681 => x"7186f40e",
  1682 => x"7e6d974d",
  1683 => x"974ca5c1",
  1684 => x"a6c8486c",
  1685 => x"c4486e58",
  1686 => x"c505a866",
  1687 => x"c048ff87",
  1688 => x"caff87e6",
  1689 => x"49a5c287",
  1690 => x"714b6c97",
  1691 => x"6b974ba3",
  1692 => x"7e6c974b",
  1693 => x"80c1486e",
  1694 => x"c758a6c8",
  1695 => x"58a6cc98",
  1696 => x"fe7c9770",
  1697 => x"487387e1",
  1698 => x"4d268ef4",
  1699 => x"4b264c26",
  1700 => x"5e0e4f26",
  1701 => x"f40e5c5b",
  1702 => x"d84c7186",
  1703 => x"ffc34a66",
  1704 => x"4ba4c29a",
  1705 => x"73496c97",
  1706 => x"517249a1",
  1707 => x"6e7e6c97",
  1708 => x"c880c148",
  1709 => x"98c758a6",
  1710 => x"7058a6cc",
  1711 => x"268ef454",
  1712 => x"264b264c",
  1713 => x"86fc1e4f",
  1714 => x"e087e4fd",
  1715 => x"c0494abf",
  1716 => x"0299c0e0",
  1717 => x"1e7287cb",
  1718 => x"49c8e8c2",
  1719 => x"c487f3fe",
  1720 => x"87fcfc86",
  1721 => x"fefc7e70",
  1722 => x"268efc87",
  1723 => x"e8c21e4f",
  1724 => x"c2fd49c8",
  1725 => x"c5ebc187",
  1726 => x"87cffc49",
  1727 => x"2687edc4",
  1728 => x"5b5e0e4f",
  1729 => x"fc0e5d5c",
  1730 => x"ff7e7186",
  1731 => x"e8c24dd4",
  1732 => x"eafc49c8",
  1733 => x"c04b7087",
  1734 => x"c204abb7",
  1735 => x"f0c387f8",
  1736 => x"87c905ab",
  1737 => x"48e4efc1",
  1738 => x"d9c278c1",
  1739 => x"abe0c387",
  1740 => x"c187c905",
  1741 => x"c148e8ef",
  1742 => x"87cac278",
  1743 => x"bfe8efc1",
  1744 => x"c287c602",
  1745 => x"c24ca3c0",
  1746 => x"c14c7387",
  1747 => x"02bfe4ef",
  1748 => x"7487e0c0",
  1749 => x"29b7c449",
  1750 => x"ecefc191",
  1751 => x"cf4a7481",
  1752 => x"c192c29a",
  1753 => x"70307248",
  1754 => x"72baff4a",
  1755 => x"70986948",
  1756 => x"7487db79",
  1757 => x"29b7c449",
  1758 => x"ecefc191",
  1759 => x"cf4a7481",
  1760 => x"c392c29a",
  1761 => x"70307248",
  1762 => x"b069484a",
  1763 => x"056e7970",
  1764 => x"ff87e7c0",
  1765 => x"e1c848d0",
  1766 => x"c17dc578",
  1767 => x"02bfe8ef",
  1768 => x"e0c387c3",
  1769 => x"e4efc17d",
  1770 => x"87c302bf",
  1771 => x"737df0c3",
  1772 => x"48d0ff7d",
  1773 => x"c078e1c8",
  1774 => x"efc178e0",
  1775 => x"78c048e8",
  1776 => x"48e4efc1",
  1777 => x"e8c278c0",
  1778 => x"f2f949c8",
  1779 => x"c04b7087",
  1780 => x"fd03abb7",
  1781 => x"48c087c8",
  1782 => x"4d268efc",
  1783 => x"4b264c26",
  1784 => x"00004f26",
  1785 => x"00000000",
  1786 => x"00000000",
  1787 => x"00000000",
  1788 => x"00000000",
  1789 => x"00000000",
  1790 => x"00000000",
  1791 => x"00000000",
  1792 => x"00000000",
  1793 => x"00000000",
  1794 => x"00000000",
  1795 => x"00000000",
  1796 => x"00000000",
  1797 => x"00000000",
  1798 => x"00000000",
  1799 => x"00000000",
  1800 => x"00000000",
  1801 => x"00000000",
  1802 => x"00000000",
  1803 => x"724ac01e",
  1804 => x"c191c449",
  1805 => x"c081ecef",
  1806 => x"d082c179",
  1807 => x"ee04aab7",
  1808 => x"0e4f2687",
  1809 => x"5d5c5b5e",
  1810 => x"f74d710e",
  1811 => x"4a7587e1",
  1812 => x"922ab7c4",
  1813 => x"82ecefc1",
  1814 => x"9ccf4c75",
  1815 => x"496a94c2",
  1816 => x"c32b744b",
  1817 => x"7448c29b",
  1818 => x"ff4c7030",
  1819 => x"714874bc",
  1820 => x"f67a7098",
  1821 => x"487387f1",
  1822 => x"4c264d26",
  1823 => x"4f264b26",
  1824 => x"48d0ff1e",
  1825 => x"7178e1c8",
  1826 => x"08d4ff48",
  1827 => x"4866c478",
  1828 => x"7808d4ff",
  1829 => x"711e4f26",
  1830 => x"4966c44a",
  1831 => x"ff49721e",
  1832 => x"d0ff87de",
  1833 => x"78e0c048",
  1834 => x"4f268efc",
  1835 => x"711e731e",
  1836 => x"4966c84b",
  1837 => x"c14a731e",
  1838 => x"ff49a2e0",
  1839 => x"8efc87d8",
  1840 => x"4f264b26",
  1841 => x"48d0ff1e",
  1842 => x"7178c9c8",
  1843 => x"08d4ff48",
  1844 => x"1e4f2678",
  1845 => x"eb494a71",
  1846 => x"48d0ff87",
  1847 => x"4f2678c8",
  1848 => x"711e731e",
  1849 => x"e0e8c24b",
  1850 => x"87c302bf",
  1851 => x"ff87ebc2",
  1852 => x"c9c848d0",
  1853 => x"c0487378",
  1854 => x"d4ffb0e0",
  1855 => x"e8c27808",
  1856 => x"78c048d4",
  1857 => x"c50266c8",
  1858 => x"49ffc387",
  1859 => x"49c087c2",
  1860 => x"59dce8c2",
  1861 => x"c60266cc",
  1862 => x"d5d5c587",
  1863 => x"cf87c44a",
  1864 => x"c24affff",
  1865 => x"c25ae0e8",
  1866 => x"c148e0e8",
  1867 => x"264b2678",
  1868 => x"5b5e0e4f",
  1869 => x"710e5d5c",
  1870 => x"dce8c24d",
  1871 => x"9d754bbf",
  1872 => x"4987cb02",
  1873 => x"f3c191c8",
  1874 => x"82714ad8",
  1875 => x"f7c187c4",
  1876 => x"4cc04ad8",
  1877 => x"99734912",
  1878 => x"bfd8e8c2",
  1879 => x"ffb87148",
  1880 => x"c17808d4",
  1881 => x"c8842bb7",
  1882 => x"e704acb7",
  1883 => x"d4e8c287",
  1884 => x"80c848bf",
  1885 => x"58d8e8c2",
  1886 => x"4c264d26",
  1887 => x"4f264b26",
  1888 => x"711e731e",
  1889 => x"9a4a134b",
  1890 => x"7287cb02",
  1891 => x"87e1fe49",
  1892 => x"059a4a13",
  1893 => x"4b2687f5",
  1894 => x"c21e4f26",
  1895 => x"49bfd4e8",
  1896 => x"48d4e8c2",
  1897 => x"c478a1c1",
  1898 => x"03a9b7c0",
  1899 => x"d4ff87db",
  1900 => x"d8e8c248",
  1901 => x"e8c278bf",
  1902 => x"c249bfd4",
  1903 => x"c148d4e8",
  1904 => x"c0c478a1",
  1905 => x"e504a9b7",
  1906 => x"48d0ff87",
  1907 => x"e8c278c8",
  1908 => x"78c048e0",
  1909 => x"00004f26",
  1910 => x"00000000",
  1911 => x"00000000",
  1912 => x"5f000000",
  1913 => x"0000005f",
  1914 => x"00030300",
  1915 => x"00000303",
  1916 => x"147f7f14",
  1917 => x"00147f7f",
  1918 => x"6b2e2400",
  1919 => x"00123a6b",
  1920 => x"18366a4c",
  1921 => x"0032566c",
  1922 => x"594f7e30",
  1923 => x"40683a77",
  1924 => x"07040000",
  1925 => x"00000003",
  1926 => x"3e1c0000",
  1927 => x"00004163",
  1928 => x"63410000",
  1929 => x"00001c3e",
  1930 => x"1c3e2a08",
  1931 => x"082a3e1c",
  1932 => x"3e080800",
  1933 => x"0008083e",
  1934 => x"e0800000",
  1935 => x"00000060",
  1936 => x"08080800",
  1937 => x"00080808",
  1938 => x"60000000",
  1939 => x"00000060",
  1940 => x"18306040",
  1941 => x"0103060c",
  1942 => x"597f3e00",
  1943 => x"003e7f4d",
  1944 => x"7f060400",
  1945 => x"0000007f",
  1946 => x"71634200",
  1947 => x"00464f59",
  1948 => x"49632200",
  1949 => x"00367f49",
  1950 => x"13161c18",
  1951 => x"00107f7f",
  1952 => x"45672700",
  1953 => x"00397d45",
  1954 => x"4b7e3c00",
  1955 => x"00307949",
  1956 => x"71010100",
  1957 => x"00070f79",
  1958 => x"497f3600",
  1959 => x"00367f49",
  1960 => x"494f0600",
  1961 => x"001e3f69",
  1962 => x"66000000",
  1963 => x"00000066",
  1964 => x"e6800000",
  1965 => x"00000066",
  1966 => x"14080800",
  1967 => x"00222214",
  1968 => x"14141400",
  1969 => x"00141414",
  1970 => x"14222200",
  1971 => x"00080814",
  1972 => x"51030200",
  1973 => x"00060f59",
  1974 => x"5d417f3e",
  1975 => x"001e1f55",
  1976 => x"097f7e00",
  1977 => x"007e7f09",
  1978 => x"497f7f00",
  1979 => x"00367f49",
  1980 => x"633e1c00",
  1981 => x"00414141",
  1982 => x"417f7f00",
  1983 => x"001c3e63",
  1984 => x"497f7f00",
  1985 => x"00414149",
  1986 => x"097f7f00",
  1987 => x"00010109",
  1988 => x"417f3e00",
  1989 => x"007a7b49",
  1990 => x"087f7f00",
  1991 => x"007f7f08",
  1992 => x"7f410000",
  1993 => x"0000417f",
  1994 => x"40602000",
  1995 => x"003f7f40",
  1996 => x"1c087f7f",
  1997 => x"00416336",
  1998 => x"407f7f00",
  1999 => x"00404040",
  2000 => x"0c067f7f",
  2001 => x"007f7f06",
  2002 => x"0c067f7f",
  2003 => x"007f7f18",
  2004 => x"417f3e00",
  2005 => x"003e7f41",
  2006 => x"097f7f00",
  2007 => x"00060f09",
  2008 => x"61417f3e",
  2009 => x"00407e7f",
  2010 => x"097f7f00",
  2011 => x"00667f19",
  2012 => x"4d6f2600",
  2013 => x"00327b59",
  2014 => x"7f010100",
  2015 => x"0001017f",
  2016 => x"407f3f00",
  2017 => x"003f7f40",
  2018 => x"703f0f00",
  2019 => x"000f3f70",
  2020 => x"18307f7f",
  2021 => x"007f7f30",
  2022 => x"1c366341",
  2023 => x"4163361c",
  2024 => x"7c060301",
  2025 => x"0103067c",
  2026 => x"4d597161",
  2027 => x"00414347",
  2028 => x"7f7f0000",
  2029 => x"00004141",
  2030 => x"0c060301",
  2031 => x"40603018",
  2032 => x"41410000",
  2033 => x"00007f7f",
  2034 => x"03060c08",
  2035 => x"00080c06",
  2036 => x"80808080",
  2037 => x"00808080",
  2038 => x"03000000",
  2039 => x"00000407",
  2040 => x"54742000",
  2041 => x"00787c54",
  2042 => x"447f7f00",
  2043 => x"00387c44",
  2044 => x"447c3800",
  2045 => x"00004444",
  2046 => x"447c3800",
  2047 => x"007f7f44",
  2048 => x"547c3800",
  2049 => x"00185c54",
  2050 => x"7f7e0400",
  2051 => x"00000505",
  2052 => x"a4bc1800",
  2053 => x"007cfca4",
  2054 => x"047f7f00",
  2055 => x"00787c04",
  2056 => x"3d000000",
  2057 => x"0000407d",
  2058 => x"80808000",
  2059 => x"00007dfd",
  2060 => x"107f7f00",
  2061 => x"00446c38",
  2062 => x"3f000000",
  2063 => x"0000407f",
  2064 => x"180c7c7c",
  2065 => x"00787c0c",
  2066 => x"047c7c00",
  2067 => x"00787c04",
  2068 => x"447c3800",
  2069 => x"00387c44",
  2070 => x"24fcfc00",
  2071 => x"00183c24",
  2072 => x"243c1800",
  2073 => x"00fcfc24",
  2074 => x"047c7c00",
  2075 => x"00080c04",
  2076 => x"545c4800",
  2077 => x"00207454",
  2078 => x"7f3f0400",
  2079 => x"00004444",
  2080 => x"407c3c00",
  2081 => x"007c7c40",
  2082 => x"603c1c00",
  2083 => x"001c3c60",
  2084 => x"30607c3c",
  2085 => x"003c7c60",
  2086 => x"10386c44",
  2087 => x"00446c38",
  2088 => x"e0bc1c00",
  2089 => x"001c3c60",
  2090 => x"74644400",
  2091 => x"00444c5c",
  2092 => x"3e080800",
  2093 => x"00414177",
  2094 => x"7f000000",
  2095 => x"0000007f",
  2096 => x"77414100",
  2097 => x"0008083e",
  2098 => x"03010102",
  2099 => x"00010202",
  2100 => x"7f7f7f7f",
  2101 => x"007f7f7f",
  2102 => x"1c1c0808",
  2103 => x"7f7f3e3e",
  2104 => x"3e3e7f7f",
  2105 => x"08081c1c",
  2106 => x"7c181000",
  2107 => x"0010187c",
  2108 => x"7c301000",
  2109 => x"0010307c",
  2110 => x"60603010",
  2111 => x"00061e78",
  2112 => x"183c6642",
  2113 => x"0042663c",
  2114 => x"c26a3878",
  2115 => x"00386cc6",
  2116 => x"60000060",
  2117 => x"00600000",
  2118 => x"5c5b5e0e",
  2119 => x"86fc0e5d",
  2120 => x"e8c27e71",
  2121 => x"c04cbfe8",
  2122 => x"c41ec04b",
  2123 => x"c402ab66",
  2124 => x"c24dc087",
  2125 => x"754dc187",
  2126 => x"ee49731e",
  2127 => x"86c887e2",
  2128 => x"ef49e0c0",
  2129 => x"a4c487eb",
  2130 => x"f0496a4a",
  2131 => x"c9f187f2",
  2132 => x"c184cc87",
  2133 => x"abb7c883",
  2134 => x"87cdff04",
  2135 => x"4d268efc",
  2136 => x"4b264c26",
  2137 => x"711e4f26",
  2138 => x"ece8c24a",
  2139 => x"ece8c25a",
  2140 => x"4978c748",
  2141 => x"2687e1fe",
  2142 => x"1e731e4f",
  2143 => x"b7c04a71",
  2144 => x"87d303aa",
  2145 => x"bff4d4c2",
  2146 => x"c187c405",
  2147 => x"c087c24b",
  2148 => x"f8d4c24b",
  2149 => x"c287c45b",
  2150 => x"fc5af8d4",
  2151 => x"f4d4c248",
  2152 => x"c14a78bf",
  2153 => x"a2c0c19a",
  2154 => x"87e7ec49",
  2155 => x"4f264b26",
  2156 => x"c44a711e",
  2157 => x"49721e66",
  2158 => x"fc87f1eb",
  2159 => x"1e4f268e",
  2160 => x"c348d4ff",
  2161 => x"d0ff78ff",
  2162 => x"78e1c048",
  2163 => x"c148d4ff",
  2164 => x"c4487178",
  2165 => x"08d4ff30",
  2166 => x"48d0ff78",
  2167 => x"2678e0c0",
  2168 => x"5b5e0e4f",
  2169 => x"f00e5d5c",
  2170 => x"48a6c886",
  2171 => x"bfec78c0",
  2172 => x"c280fc7e",
  2173 => x"78bfe8e8",
  2174 => x"bff0e8c2",
  2175 => x"4cbfe84d",
  2176 => x"bff4d4c2",
  2177 => x"87f9e349",
  2178 => x"f6e849c7",
  2179 => x"c2497087",
  2180 => x"87cf0599",
  2181 => x"bfecd4c2",
  2182 => x"6eb9ff49",
  2183 => x"0299c199",
  2184 => x"cb87c0c2",
  2185 => x"cfcc49ee",
  2186 => x"58a6d087",
  2187 => x"d2e849c7",
  2188 => x"05987087",
  2189 => x"496e87c8",
  2190 => x"c10299c1",
  2191 => x"66cc87c2",
  2192 => x"7ebfec4b",
  2193 => x"bff4d4c2",
  2194 => x"87f5e249",
  2195 => x"f3cb4973",
  2196 => x"02987087",
  2197 => x"d4c287d7",
  2198 => x"c149bfd4",
  2199 => x"d8d4c2b9",
  2200 => x"dafd7159",
  2201 => x"49eecb87",
  2202 => x"7087cdcb",
  2203 => x"e749c74b",
  2204 => x"987087d1",
  2205 => x"87c9ff05",
  2206 => x"99c1496e",
  2207 => x"87c1ff05",
  2208 => x"bff4d4c2",
  2209 => x"c2bac14a",
  2210 => x"fc5af8d4",
  2211 => x"c10a7a0a",
  2212 => x"a2c0c19a",
  2213 => x"87fbe849",
  2214 => x"e649dac1",
  2215 => x"a6c887e5",
  2216 => x"c278c148",
  2217 => x"6e48ecd4",
  2218 => x"f4d4c278",
  2219 => x"c7c105bf",
  2220 => x"c0c0c887",
  2221 => x"e0d5c24b",
  2222 => x"49154d7e",
  2223 => x"87c3e649",
  2224 => x"c0029870",
  2225 => x"b47387c2",
  2226 => x"052bb7c1",
  2227 => x"7487ebff",
  2228 => x"99ffc349",
  2229 => x"49c01e71",
  2230 => x"7487d5fb",
  2231 => x"29b7c849",
  2232 => x"49c11e71",
  2233 => x"c887c9fb",
  2234 => x"49fdc386",
  2235 => x"c387d4e5",
  2236 => x"cee549fa",
  2237 => x"87d1c887",
  2238 => x"ffc34974",
  2239 => x"2cb7c899",
  2240 => x"9c74b471",
  2241 => x"ff87df02",
  2242 => x"497ebfc8",
  2243 => x"bff0d4c2",
  2244 => x"a9e0c289",
  2245 => x"87c5c003",
  2246 => x"cfc04cc0",
  2247 => x"f0d4c287",
  2248 => x"c0786e48",
  2249 => x"d4c287c6",
  2250 => x"78c048f0",
  2251 => x"99c84974",
  2252 => x"87cec005",
  2253 => x"e449f5c3",
  2254 => x"497087c9",
  2255 => x"c00299c2",
  2256 => x"e8c287ea",
  2257 => x"c002bfec",
  2258 => x"c14887ca",
  2259 => x"f0e8c288",
  2260 => x"87d3c058",
  2261 => x"c14866c4",
  2262 => x"7e7080e0",
  2263 => x"c002bf6e",
  2264 => x"ff4b87c5",
  2265 => x"c80f7349",
  2266 => x"78c148a6",
  2267 => x"99c44974",
  2268 => x"87cec005",
  2269 => x"e349f2c3",
  2270 => x"497087c9",
  2271 => x"c00299c2",
  2272 => x"e8c287f0",
  2273 => x"487ebfec",
  2274 => x"03a8b7c7",
  2275 => x"6e87cbc0",
  2276 => x"c280c148",
  2277 => x"c058f0e8",
  2278 => x"66c487d3",
  2279 => x"80e0c148",
  2280 => x"bf6e7e70",
  2281 => x"87c5c002",
  2282 => x"7349fe4b",
  2283 => x"48a6c80f",
  2284 => x"fdc378c1",
  2285 => x"87cbe249",
  2286 => x"99c24970",
  2287 => x"87e6c002",
  2288 => x"bfece8c2",
  2289 => x"87c9c002",
  2290 => x"48ece8c2",
  2291 => x"d0c078c0",
  2292 => x"4a66c487",
  2293 => x"6a82e0c1",
  2294 => x"87c5c002",
  2295 => x"7349fd4b",
  2296 => x"48a6c80f",
  2297 => x"fac378c1",
  2298 => x"87d7e149",
  2299 => x"99c24970",
  2300 => x"87edc002",
  2301 => x"bfece8c2",
  2302 => x"a8b7c748",
  2303 => x"87c9c003",
  2304 => x"48ece8c2",
  2305 => x"d3c078c7",
  2306 => x"4866c487",
  2307 => x"7080e0c1",
  2308 => x"02bf6e7e",
  2309 => x"4b87c5c0",
  2310 => x"0f7349fc",
  2311 => x"c148a6c8",
  2312 => x"c3487478",
  2313 => x"7e7098f0",
  2314 => x"c0059848",
  2315 => x"dac187ce",
  2316 => x"87cfe049",
  2317 => x"99c24970",
  2318 => x"87d0c202",
  2319 => x"c349eecb",
  2320 => x"a6d087f6",
  2321 => x"e4e8c258",
  2322 => x"c250c048",
  2323 => x"bf97e4e8",
  2324 => x"87d8c105",
  2325 => x"cdc0056e",
  2326 => x"49dac187",
  2327 => x"87e3dfff",
  2328 => x"c1029870",
  2329 => x"bfe887c6",
  2330 => x"ffc3494b",
  2331 => x"2bb7c899",
  2332 => x"d4c2b371",
  2333 => x"ff49bff4",
  2334 => x"cc87c6da",
  2335 => x"c3c34966",
  2336 => x"02987087",
  2337 => x"c287c6c0",
  2338 => x"c148e4e8",
  2339 => x"e4e8c250",
  2340 => x"c005bf97",
  2341 => x"497387d6",
  2342 => x"0599f0c3",
  2343 => x"c187c7ff",
  2344 => x"deff49da",
  2345 => x"987087dd",
  2346 => x"87fafe05",
  2347 => x"c248a6cc",
  2348 => x"78bfece8",
  2349 => x"cc4966cc",
  2350 => x"4866c491",
  2351 => x"7e708071",
  2352 => x"c002bf6e",
  2353 => x"cc4b87c6",
  2354 => x"0f734966",
  2355 => x"c0029d75",
  2356 => x"026d87e9",
  2357 => x"6d87e4c0",
  2358 => x"e6ddff49",
  2359 => x"c1497087",
  2360 => x"cbc00299",
  2361 => x"4ba5c487",
  2362 => x"bfece8c2",
  2363 => x"0f4b6b49",
  2364 => x"c00285c8",
  2365 => x"056d87c5",
  2366 => x"c887dcff",
  2367 => x"c8c00266",
  2368 => x"ece8c287",
  2369 => x"cff049bf",
  2370 => x"268ef087",
  2371 => x"264c264d",
  2372 => x"004f264b",
  2373 => x"00000000",
  2374 => x"00000010",
  2375 => x"14111258",
  2376 => x"231c1b1d",
  2377 => x"9491595a",
  2378 => x"f4ebf2f5",
  2379 => x"00000000",
  2380 => x"00000000",
  2381 => x"00000000",
  2382 => x"ff4a711e",
  2383 => x"7249bfc8",
  2384 => x"4f2648a1",
  2385 => x"bfc8ff1e",
  2386 => x"c0c0fe89",
  2387 => x"a9c0c0c0",
  2388 => x"c087c401",
  2389 => x"c187c24a",
  2390 => x"2648724a",
  2391 => x"0000004f",
  2392 => x"11141258",
  2393 => x"231c1b1d",
  2394 => x"9194595a",
  2395 => x"f4ebf2f5",
  2396 => x"00002574",
  2397 => x"4f545541",
  2398 => x"544f4f42",
  2399 => x"17004247",
  2400 => x"1700001a",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
