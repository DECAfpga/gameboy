library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"f8e6c287",
    12 => x"48c0c84e",
    13 => x"d5c128c2",
    14 => x"ead6e5ea",
    15 => x"c1467149",
    16 => x"87f90188",
    17 => x"49f8e6c2",
    18 => x"48f4d3c2",
    19 => x"0389d089",
    20 => x"404040c0",
    21 => x"d087f640",
    22 => x"50c00581",
    23 => x"f90589c1",
    24 => x"f3d3c287",
    25 => x"efd3c24d",
    26 => x"02ad744c",
    27 => x"0f2487c4",
    28 => x"e0c187f7",
    29 => x"d3c287ef",
    30 => x"d3c24df3",
    31 => x"ad744cf3",
    32 => x"c487c602",
    33 => x"f50f6c8c",
    34 => x"87fd0087",
    35 => x"7186fc1e",
    36 => x"49c0ff4a",
    37 => x"c0c44869",
    38 => x"487e7098",
    39 => x"87f40298",
    40 => x"fc487972",
    41 => x"0e4f268e",
    42 => x"0e5c5b5e",
    43 => x"4cc04b71",
    44 => x"029a4a13",
    45 => x"497287cd",
    46 => x"c187d1ff",
    47 => x"9a4a1384",
    48 => x"7487f305",
    49 => x"264c2648",
    50 => x"1e4f264b",
    51 => x"1e731e72",
    52 => x"02114812",
    53 => x"c34b87ca",
    54 => x"739b98df",
    55 => x"87f00288",
    56 => x"4a264b26",
    57 => x"731e4f26",
    58 => x"c11e721e",
    59 => x"87ca048b",
    60 => x"02114812",
    61 => x"028887c4",
    62 => x"4a2687f1",
    63 => x"4f264b26",
    64 => x"731e741e",
    65 => x"c11e721e",
    66 => x"87cf048b",
    67 => x"02114812",
    68 => x"df4c87c9",
    69 => x"88749c98",
    70 => x"2687ec02",
    71 => x"264b264a",
    72 => x"1e4f264c",
    73 => x"73814873",
    74 => x"87c502a9",
    75 => x"f6055312",
    76 => x"0e4f2687",
    77 => x"0e5c5b5e",
    78 => x"d4ff4a71",
    79 => x"4b66cc4c",
    80 => x"718bc149",
    81 => x"87ce0299",
    82 => x"6c7cffc3",
    83 => x"c1497352",
    84 => x"0599718b",
    85 => x"4c2687f2",
    86 => x"4f264b26",
    87 => x"ff1e731e",
    88 => x"ffc34bd4",
    89 => x"c34a6b7b",
    90 => x"496b7bff",
    91 => x"b17232c8",
    92 => x"6b7bffc3",
    93 => x"7131c84a",
    94 => x"7bffc3b2",
    95 => x"32c8496b",
    96 => x"4871b172",
    97 => x"4f264b26",
    98 => x"5c5b5e0e",
    99 => x"4d710e5d",
   100 => x"754cd4ff",
   101 => x"98ffc348",
   102 => x"d3c27c70",
   103 => x"c805bff4",
   104 => x"4866d087",
   105 => x"a6d430c9",
   106 => x"4966d058",
   107 => x"487129d8",
   108 => x"7098ffc3",
   109 => x"4966d07c",
   110 => x"487129d0",
   111 => x"7098ffc3",
   112 => x"4966d07c",
   113 => x"487129c8",
   114 => x"7098ffc3",
   115 => x"4866d07c",
   116 => x"7098ffc3",
   117 => x"d049757c",
   118 => x"c3487129",
   119 => x"7c7098ff",
   120 => x"f0c94b6c",
   121 => x"ffc34aff",
   122 => x"87cf05ab",
   123 => x"6c7c7149",
   124 => x"028ac14b",
   125 => x"ab7187c5",
   126 => x"7387f202",
   127 => x"264d2648",
   128 => x"264b264c",
   129 => x"49c01e4f",
   130 => x"c348d4ff",
   131 => x"81c178ff",
   132 => x"a9b7c8c3",
   133 => x"2687f104",
   134 => x"5b5e0e4f",
   135 => x"c00e5d5c",
   136 => x"f7c1f0ff",
   137 => x"c0c0c14d",
   138 => x"4bc0c0c0",
   139 => x"c487d6ff",
   140 => x"c04cdff8",
   141 => x"fd49751e",
   142 => x"86c487ce",
   143 => x"c005a8c1",
   144 => x"d4ff87e5",
   145 => x"78ffc348",
   146 => x"e1c01e73",
   147 => x"49e9c1f0",
   148 => x"c487f5fc",
   149 => x"05987086",
   150 => x"d4ff87ca",
   151 => x"78ffc348",
   152 => x"87cb48c1",
   153 => x"c187defe",
   154 => x"c6ff058c",
   155 => x"2648c087",
   156 => x"264c264d",
   157 => x"0e4f264b",
   158 => x"0e5c5b5e",
   159 => x"c1f0ffc0",
   160 => x"d4ff4cc1",
   161 => x"78ffc348",
   162 => x"f849fcca",
   163 => x"4bd387d9",
   164 => x"49741ec0",
   165 => x"c487f1fb",
   166 => x"05987086",
   167 => x"d4ff87ca",
   168 => x"78ffc348",
   169 => x"87cb48c1",
   170 => x"c187dafd",
   171 => x"dfff058b",
   172 => x"2648c087",
   173 => x"264b264c",
   174 => x"0000004f",
   175 => x"00444d43",
   176 => x"43484453",
   177 => x"69616620",
   178 => x"000a216c",
   179 => x"52524549",
   180 => x"00000000",
   181 => x"00495053",
   182 => x"74697257",
   183 => x"61662065",
   184 => x"64656c69",
   185 => x"5e0e000a",
   186 => x"0e5d5c5b",
   187 => x"ff4dffc3",
   188 => x"d0fc4bd4",
   189 => x"1eeac687",
   190 => x"c1f0e1c0",
   191 => x"c7fa49c8",
   192 => x"c186c487",
   193 => x"87c802a8",
   194 => x"c087ecfd",
   195 => x"87e8c148",
   196 => x"7087c9f9",
   197 => x"ffffcf49",
   198 => x"a9eac699",
   199 => x"fd87c802",
   200 => x"48c087d5",
   201 => x"7587d1c1",
   202 => x"4cf1c07b",
   203 => x"7087eafb",
   204 => x"ecc00298",
   205 => x"c01ec087",
   206 => x"fac1f0ff",
   207 => x"87c8f949",
   208 => x"987086c4",
   209 => x"7587da05",
   210 => x"75496b7b",
   211 => x"757b757b",
   212 => x"c17b757b",
   213 => x"c40299c0",
   214 => x"db48c187",
   215 => x"d748c087",
   216 => x"05acc287",
   217 => x"c0cb87ca",
   218 => x"87fbf449",
   219 => x"87c848c0",
   220 => x"fe058cc1",
   221 => x"48c087f6",
   222 => x"4c264d26",
   223 => x"4f264b26",
   224 => x"5c5b5e0e",
   225 => x"d0ff0e5d",
   226 => x"d0e5c04d",
   227 => x"c24cc0c1",
   228 => x"c148f4d3",
   229 => x"49d4cb78",
   230 => x"c787ccf4",
   231 => x"f97dc24b",
   232 => x"7dc387e3",
   233 => x"49741ec0",
   234 => x"c487ddf7",
   235 => x"05a8c186",
   236 => x"c24b87c1",
   237 => x"87cb05ab",
   238 => x"f349cccb",
   239 => x"48c087e9",
   240 => x"c187f6c0",
   241 => x"d4ff058b",
   242 => x"87dafc87",
   243 => x"58f8d3c2",
   244 => x"cd059870",
   245 => x"c01ec187",
   246 => x"d0c1f0ff",
   247 => x"87e8f649",
   248 => x"d4ff86c4",
   249 => x"78ffc348",
   250 => x"c287c3c3",
   251 => x"c258fcd3",
   252 => x"48d4ff7d",
   253 => x"c178ffc3",
   254 => x"264d2648",
   255 => x"264b264c",
   256 => x"5b5e0e4f",
   257 => x"fc0e5d5c",
   258 => x"ff4b7186",
   259 => x"7ec04cd4",
   260 => x"dfcdeec5",
   261 => x"7cffc34a",
   262 => x"fec3486c",
   263 => x"f8c005a8",
   264 => x"734d7487",
   265 => x"87cc029b",
   266 => x"731e66d4",
   267 => x"87c3f449",
   268 => x"87d486c4",
   269 => x"c448d0ff",
   270 => x"66d478d1",
   271 => x"7dffc34a",
   272 => x"f8058ac1",
   273 => x"5aa6d887",
   274 => x"7c7cffc3",
   275 => x"c5059b73",
   276 => x"48d0ff87",
   277 => x"4ac178d0",
   278 => x"058ac17e",
   279 => x"6e87f6fe",
   280 => x"268efc48",
   281 => x"264c264d",
   282 => x"1e4f264b",
   283 => x"4a711e73",
   284 => x"d4ff4bc0",
   285 => x"78ffc348",
   286 => x"c448d0ff",
   287 => x"d4ff78c3",
   288 => x"78ffc348",
   289 => x"ffc01e72",
   290 => x"49d1c1f0",
   291 => x"c487f9f3",
   292 => x"05987086",
   293 => x"c0c887d2",
   294 => x"4966cc1e",
   295 => x"c487e2fd",
   296 => x"ff4b7086",
   297 => x"78c248d0",
   298 => x"4b264873",
   299 => x"5e0e4f26",
   300 => x"0e5d5c5b",
   301 => x"ffc01ec0",
   302 => x"49c9c1f0",
   303 => x"d287c9f3",
   304 => x"c4d4c21e",
   305 => x"87f9fc49",
   306 => x"4cc086c8",
   307 => x"b7d284c1",
   308 => x"87f804ac",
   309 => x"97c4d4c2",
   310 => x"c0c349bf",
   311 => x"a9c0c199",
   312 => x"87e7c005",
   313 => x"97cbd4c2",
   314 => x"31d049bf",
   315 => x"97ccd4c2",
   316 => x"32c84abf",
   317 => x"d4c2b172",
   318 => x"4abf97cd",
   319 => x"cf4c71b1",
   320 => x"9cffffff",
   321 => x"34ca84c1",
   322 => x"c287e7c1",
   323 => x"bf97cdd4",
   324 => x"c631c149",
   325 => x"ced4c299",
   326 => x"c74abf97",
   327 => x"b1722ab7",
   328 => x"97c9d4c2",
   329 => x"cf4d4abf",
   330 => x"cad4c29d",
   331 => x"c34abf97",
   332 => x"c232ca9a",
   333 => x"bf97cbd4",
   334 => x"7333c24b",
   335 => x"ccd4c2b2",
   336 => x"c34bbf97",
   337 => x"b7c69bc0",
   338 => x"c2b2732b",
   339 => x"7148c181",
   340 => x"c1497030",
   341 => x"70307548",
   342 => x"c14c724d",
   343 => x"c8947184",
   344 => x"06adb7c0",
   345 => x"34c187cc",
   346 => x"c0c82db7",
   347 => x"ff01adb7",
   348 => x"487487f4",
   349 => x"4c264d26",
   350 => x"4f264b26",
   351 => x"5c5b5e0e",
   352 => x"86fc0e5d",
   353 => x"48ecdcc2",
   354 => x"d4c278c0",
   355 => x"49c01ee4",
   356 => x"c487d8fb",
   357 => x"05987086",
   358 => x"48c087c5",
   359 => x"c087d1c9",
   360 => x"e8e1c24d",
   361 => x"c278c148",
   362 => x"c04adad5",
   363 => x"c849c8e0",
   364 => x"87f2ec4b",
   365 => x"c6059870",
   366 => x"e8e1c287",
   367 => x"c278c048",
   368 => x"c04af6d5",
   369 => x"c849d4e0",
   370 => x"87daec4b",
   371 => x"c6059870",
   372 => x"e8e1c287",
   373 => x"c278c048",
   374 => x"02bfe8e1",
   375 => x"c287fdc0",
   376 => x"4dbfeadb",
   377 => x"9fe2dcc2",
   378 => x"c5487ebf",
   379 => x"05a8ead6",
   380 => x"dbc287c7",
   381 => x"ce4dbfea",
   382 => x"ca486e87",
   383 => x"02a8d5e9",
   384 => x"48c087c5",
   385 => x"c287e9c7",
   386 => x"751ee4d4",
   387 => x"87dbf949",
   388 => x"987086c4",
   389 => x"c087c505",
   390 => x"87d4c748",
   391 => x"4af6d5c2",
   392 => x"49e0e0c0",
   393 => x"fdea4bc8",
   394 => x"05987087",
   395 => x"dcc287c8",
   396 => x"78c148ec",
   397 => x"d5c287d8",
   398 => x"e0c04ada",
   399 => x"4bc849ec",
   400 => x"7087e3ea",
   401 => x"c5c00298",
   402 => x"c648c087",
   403 => x"dcc287e2",
   404 => x"49bf97e2",
   405 => x"05a9d5c1",
   406 => x"c287cdc0",
   407 => x"bf97e3dc",
   408 => x"a9eac249",
   409 => x"87c5c002",
   410 => x"c3c648c0",
   411 => x"e4d4c287",
   412 => x"487ebf97",
   413 => x"02a8e9c3",
   414 => x"6e87cec0",
   415 => x"a8ebc348",
   416 => x"87c5c002",
   417 => x"e7c548c0",
   418 => x"efd4c287",
   419 => x"9949bf97",
   420 => x"87ccc005",
   421 => x"97f0d4c2",
   422 => x"a9c249bf",
   423 => x"87c5c002",
   424 => x"cbc548c0",
   425 => x"f1d4c287",
   426 => x"c248bf97",
   427 => x"7058e8dc",
   428 => x"88c1484c",
   429 => x"58ecdcc2",
   430 => x"97f2d4c2",
   431 => x"817549bf",
   432 => x"97f3d4c2",
   433 => x"32c84abf",
   434 => x"c27ea172",
   435 => x"6e48c4e1",
   436 => x"f4d4c278",
   437 => x"c248bf97",
   438 => x"c258dce1",
   439 => x"02bfecdc",
   440 => x"c287d2c2",
   441 => x"df4af6d5",
   442 => x"4bc849fc",
   443 => x"7087f7e7",
   444 => x"c5c00298",
   445 => x"c348c087",
   446 => x"dcc287f6",
   447 => x"c24cbfe4",
   448 => x"c25cd8e1",
   449 => x"bf97c9d5",
   450 => x"c231c849",
   451 => x"bf97c8d5",
   452 => x"c249a14a",
   453 => x"bf97cad5",
   454 => x"7232d04a",
   455 => x"d5c249a1",
   456 => x"4abf97cb",
   457 => x"a17232d8",
   458 => x"e0e1c249",
   459 => x"d8e1c259",
   460 => x"e1c291bf",
   461 => x"c281bfc4",
   462 => x"c259cce1",
   463 => x"bf97d1d5",
   464 => x"c232c84a",
   465 => x"bf97d0d5",
   466 => x"c24aa24b",
   467 => x"bf97d2d5",
   468 => x"7333d04b",
   469 => x"d5c24aa2",
   470 => x"4bbf97d3",
   471 => x"33d89bcf",
   472 => x"c24aa273",
   473 => x"c25ad0e1",
   474 => x"c292748a",
   475 => x"7248d0e1",
   476 => x"c7c178a1",
   477 => x"f6d4c287",
   478 => x"c849bf97",
   479 => x"f5d4c231",
   480 => x"a14abf97",
   481 => x"c731c549",
   482 => x"29c981ff",
   483 => x"59d8e1c2",
   484 => x"97fbd4c2",
   485 => x"32c84abf",
   486 => x"97fad4c2",
   487 => x"4aa24bbf",
   488 => x"5ae0e1c2",
   489 => x"bfd8e1c2",
   490 => x"c2826e92",
   491 => x"c25ad4e1",
   492 => x"c048cce1",
   493 => x"c8e1c278",
   494 => x"78a17248",
   495 => x"48e0e1c2",
   496 => x"bfcce1c2",
   497 => x"e4e1c278",
   498 => x"d0e1c248",
   499 => x"dcc278bf",
   500 => x"c002bfec",
   501 => x"487487c9",
   502 => x"7e7030c4",
   503 => x"c287c9c0",
   504 => x"48bfd4e1",
   505 => x"7e7030c4",
   506 => x"48f0dcc2",
   507 => x"48c1786e",
   508 => x"4d268efc",
   509 => x"4b264c26",
   510 => x"00004f26",
   511 => x"33544146",
   512 => x"20202032",
   513 => x"00000000",
   514 => x"31544146",
   515 => x"20202036",
   516 => x"00000000",
   517 => x"33544146",
   518 => x"20202032",
   519 => x"00000000",
   520 => x"33544146",
   521 => x"20202032",
   522 => x"00000000",
   523 => x"31544146",
   524 => x"20202036",
   525 => x"5b5e0e00",
   526 => x"710e5d5c",
   527 => x"ecdcc24a",
   528 => x"87cb02bf",
   529 => x"2bc74b72",
   530 => x"ffc14d72",
   531 => x"7287c99d",
   532 => x"722bc84b",
   533 => x"9dffc34d",
   534 => x"bfc4e1c2",
   535 => x"c0f2c083",
   536 => x"d902abbf",
   537 => x"c4f2c087",
   538 => x"e4d4c25b",
   539 => x"ef49731e",
   540 => x"86c487f9",
   541 => x"c5059870",
   542 => x"c048c087",
   543 => x"dcc287e6",
   544 => x"d202bfec",
   545 => x"c4497587",
   546 => x"e4d4c291",
   547 => x"cf4c6981",
   548 => x"ffffffff",
   549 => x"7587cb9c",
   550 => x"c291c249",
   551 => x"9f81e4d4",
   552 => x"48744c69",
   553 => x"4c264d26",
   554 => x"4f264b26",
   555 => x"5c5b5e0e",
   556 => x"86f40e5d",
   557 => x"c859a6cc",
   558 => x"80c84866",
   559 => x"c0487e70",
   560 => x"49c11e78",
   561 => x"87c1c749",
   562 => x"4c7086c4",
   563 => x"fbc0029c",
   564 => x"f4dcc287",
   565 => x"4966dc4a",
   566 => x"87efdfff",
   567 => x"c0029870",
   568 => x"4a7487ea",
   569 => x"cb4966dc",
   570 => x"87d4e04b",
   571 => x"db029870",
   572 => x"741ec087",
   573 => x"87c4029c",
   574 => x"87c24dc0",
   575 => x"49754dc1",
   576 => x"c487c6c6",
   577 => x"9c4c7086",
   578 => x"87c5ff05",
   579 => x"c1029c74",
   580 => x"a4dc87d7",
   581 => x"69486e49",
   582 => x"49a4da78",
   583 => x"c44866c8",
   584 => x"58a6c880",
   585 => x"c448699f",
   586 => x"c2780866",
   587 => x"02bfecdc",
   588 => x"a4d487d2",
   589 => x"49699f49",
   590 => x"99ffffc0",
   591 => x"30d04871",
   592 => x"87c27e70",
   593 => x"486e7ec0",
   594 => x"80bf66c4",
   595 => x"780866c4",
   596 => x"c04866c8",
   597 => x"4966c878",
   598 => x"66c481cc",
   599 => x"66c879bf",
   600 => x"c081d049",
   601 => x"c248c179",
   602 => x"f448c087",
   603 => x"264d268e",
   604 => x"264b264c",
   605 => x"5b5e0e4f",
   606 => x"710e5d5c",
   607 => x"4d66d04c",
   608 => x"72496c4a",
   609 => x"c2b94da1",
   610 => x"4abfe8dc",
   611 => x"9972baff",
   612 => x"c0029971",
   613 => x"a4c487e4",
   614 => x"fa496b4b",
   615 => x"7b7087d7",
   616 => x"bfe4dcc2",
   617 => x"71816c49",
   618 => x"c2b9757c",
   619 => x"4abfe8dc",
   620 => x"9972baff",
   621 => x"ff059971",
   622 => x"7c7587dc",
   623 => x"4c264d26",
   624 => x"4f264b26",
   625 => x"711e731e",
   626 => x"c8e1c24b",
   627 => x"a3c449bf",
   628 => x"c24a6a4a",
   629 => x"e4dcc28a",
   630 => x"a17292bf",
   631 => x"e8dcc249",
   632 => x"9a6b4abf",
   633 => x"c049a172",
   634 => x"c859c4f2",
   635 => x"e9711e66",
   636 => x"86c487f9",
   637 => x"c4059870",
   638 => x"c248c087",
   639 => x"2648c187",
   640 => x"0e4f264b",
   641 => x"0e5c5b5e",
   642 => x"4bc04a71",
   643 => x"c0029a72",
   644 => x"a2da87e0",
   645 => x"4b699f49",
   646 => x"bfecdcc2",
   647 => x"d487cf02",
   648 => x"699f49a2",
   649 => x"ffc04c49",
   650 => x"34d09cff",
   651 => x"4cc087c2",
   652 => x"9b73b374",
   653 => x"4a87df02",
   654 => x"dcc28ac2",
   655 => x"9249bfe4",
   656 => x"bfc8e1c2",
   657 => x"c2807248",
   658 => x"7158e8e1",
   659 => x"c230c448",
   660 => x"c058f4dc",
   661 => x"e1c287e9",
   662 => x"c24bbfcc",
   663 => x"c248e4e1",
   664 => x"78bfd0e1",
   665 => x"bfecdcc2",
   666 => x"c287c902",
   667 => x"49bfe4dc",
   668 => x"87c731c4",
   669 => x"bfd4e1c2",
   670 => x"c231c449",
   671 => x"c259f4dc",
   672 => x"265be4e1",
   673 => x"264b264c",
   674 => x"5b5e0e4f",
   675 => x"f00e5d5c",
   676 => x"59a6c886",
   677 => x"ffffffcf",
   678 => x"7ec04cf8",
   679 => x"d80266c4",
   680 => x"e0d4c287",
   681 => x"c278c048",
   682 => x"c248d8d4",
   683 => x"78bfe4e1",
   684 => x"48dcd4c2",
   685 => x"bfe0e1c2",
   686 => x"c1ddc278",
   687 => x"c250c048",
   688 => x"49bff0dc",
   689 => x"bfe0d4c2",
   690 => x"03aa714a",
   691 => x"7287cbc4",
   692 => x"0599cf49",
   693 => x"c087e9c0",
   694 => x"c248c0f2",
   695 => x"78bfd8d4",
   696 => x"1ee4d4c2",
   697 => x"bfd8d4c2",
   698 => x"d8d4c249",
   699 => x"78a1c148",
   700 => x"87f7e571",
   701 => x"f1c086c4",
   702 => x"d4c248fc",
   703 => x"87cc78e4",
   704 => x"bffcf1c0",
   705 => x"80e0c048",
   706 => x"58c0f2c0",
   707 => x"bfe0d4c2",
   708 => x"c280c148",
   709 => x"2758e4d4",
   710 => x"00000c7c",
   711 => x"4dbf97bf",
   712 => x"e5c2029d",
   713 => x"ade5c387",
   714 => x"87dec202",
   715 => x"bffcf1c0",
   716 => x"49a3cb4b",
   717 => x"accf4c11",
   718 => x"87d2c105",
   719 => x"99df4975",
   720 => x"91cd89c1",
   721 => x"81f4dcc2",
   722 => x"124aa3c1",
   723 => x"4aa3c351",
   724 => x"a3c55112",
   725 => x"c751124a",
   726 => x"51124aa3",
   727 => x"124aa3c9",
   728 => x"4aa3ce51",
   729 => x"a3d05112",
   730 => x"d251124a",
   731 => x"51124aa3",
   732 => x"124aa3d4",
   733 => x"4aa3d651",
   734 => x"a3d85112",
   735 => x"dc51124a",
   736 => x"51124aa3",
   737 => x"124aa3de",
   738 => x"c07ec151",
   739 => x"497487fc",
   740 => x"c00599c8",
   741 => x"497487ed",
   742 => x"d30599d0",
   743 => x"66e0c087",
   744 => x"87ccc002",
   745 => x"e0c04973",
   746 => x"98700f66",
   747 => x"87d3c002",
   748 => x"c6c0056e",
   749 => x"f4dcc287",
   750 => x"c050c048",
   751 => x"48bffcf1",
   752 => x"c287e9c2",
   753 => x"c048c1dd",
   754 => x"dcc27e50",
   755 => x"c249bff0",
   756 => x"4abfe0d4",
   757 => x"fb04aa71",
   758 => x"ffcf87f5",
   759 => x"4cf8ffff",
   760 => x"bfe4e1c2",
   761 => x"87c8c005",
   762 => x"bfecdcc2",
   763 => x"87fac102",
   764 => x"bfdcd4c2",
   765 => x"87fdf049",
   766 => x"58e0d4c2",
   767 => x"c248a6c4",
   768 => x"78bfdcd4",
   769 => x"bfecdcc2",
   770 => x"87dbc002",
   771 => x"744966c4",
   772 => x"02a97499",
   773 => x"c887c8c0",
   774 => x"78c048a6",
   775 => x"c887e7c0",
   776 => x"78c148a6",
   777 => x"c487dfc0",
   778 => x"ffcf4966",
   779 => x"02a999f8",
   780 => x"cc87c8c0",
   781 => x"78c048a6",
   782 => x"cc87c5c0",
   783 => x"78c148a6",
   784 => x"cc48a6c8",
   785 => x"66c87866",
   786 => x"87dec005",
   787 => x"c24966c4",
   788 => x"e4dcc289",
   789 => x"e1c291bf",
   790 => x"7148bfc8",
   791 => x"dcd4c280",
   792 => x"e0d4c258",
   793 => x"f978c048",
   794 => x"48c087d5",
   795 => x"ffffffcf",
   796 => x"8ef04cf8",
   797 => x"4c264d26",
   798 => x"4f264b26",
   799 => x"00000000",
   800 => x"ffffffff",
   801 => x"48d4ff1e",
   802 => x"6878ffc3",
   803 => x"1e4f2648",
   804 => x"c348d4ff",
   805 => x"d0ff78ff",
   806 => x"78e1c048",
   807 => x"d448d4ff",
   808 => x"1e4f2678",
   809 => x"c048d0ff",
   810 => x"4f2678e0",
   811 => x"87d4ff1e",
   812 => x"02994970",
   813 => x"fbc087c6",
   814 => x"87f105a9",
   815 => x"4f264871",
   816 => x"5c5b5e0e",
   817 => x"c04b710e",
   818 => x"87f8fe4c",
   819 => x"02994970",
   820 => x"c087f9c0",
   821 => x"c002a9ec",
   822 => x"fbc087f2",
   823 => x"ebc002a9",
   824 => x"b766cc87",
   825 => x"87c703ac",
   826 => x"c20266d0",
   827 => x"71537187",
   828 => x"87c20299",
   829 => x"cbfe84c1",
   830 => x"99497087",
   831 => x"c087cd02",
   832 => x"c702a9ec",
   833 => x"a9fbc087",
   834 => x"87d5ff05",
   835 => x"c30266d0",
   836 => x"7b97c087",
   837 => x"05a9ecc0",
   838 => x"4a7487c4",
   839 => x"4a7487c5",
   840 => x"728a0ac0",
   841 => x"264c2648",
   842 => x"1e4f264b",
   843 => x"7087d5fd",
   844 => x"f0c04a49",
   845 => x"87c904aa",
   846 => x"01aaf9c0",
   847 => x"f0c087c3",
   848 => x"aac1c18a",
   849 => x"c187c904",
   850 => x"c301aada",
   851 => x"8af7c087",
   852 => x"4f264872",
   853 => x"5c5b5e0e",
   854 => x"86f80e5d",
   855 => x"7ec04c71",
   856 => x"c087ecfc",
   857 => x"f4f7c04b",
   858 => x"c049bf97",
   859 => x"87cf04a9",
   860 => x"c187f9fc",
   861 => x"f4f7c083",
   862 => x"ab49bf97",
   863 => x"c087f106",
   864 => x"bf97f4f7",
   865 => x"fb87cf02",
   866 => x"497087fa",
   867 => x"87c60299",
   868 => x"05a9ecc0",
   869 => x"4bc087f1",
   870 => x"7087e9fb",
   871 => x"87e4fb4d",
   872 => x"fb58a6c8",
   873 => x"4a7087de",
   874 => x"a4c883c1",
   875 => x"49699749",
   876 => x"87da05ad",
   877 => x"9749a4c9",
   878 => x"66c44969",
   879 => x"87ce05a9",
   880 => x"9749a4ca",
   881 => x"05aa4969",
   882 => x"7ec187c4",
   883 => x"ecc087d0",
   884 => x"87c602ad",
   885 => x"05adfbc0",
   886 => x"4bc087c4",
   887 => x"026e7ec1",
   888 => x"fa87f5fe",
   889 => x"487387fd",
   890 => x"4d268ef8",
   891 => x"4b264c26",
   892 => x"00004f26",
   893 => x"1e731e00",
   894 => x"c84bd4ff",
   895 => x"d0ff4a66",
   896 => x"78c5c848",
   897 => x"c148d4ff",
   898 => x"7b1178d4",
   899 => x"f9058ac1",
   900 => x"48d0ff87",
   901 => x"4b2678c4",
   902 => x"5e0e4f26",
   903 => x"0e5d5c5b",
   904 => x"7e7186f8",
   905 => x"e1c21e6e",
   906 => x"ffe949f8",
   907 => x"7086c487",
   908 => x"e4c40298",
   909 => x"e0e4c187",
   910 => x"496e4cbf",
   911 => x"c887d5fc",
   912 => x"987058a6",
   913 => x"c487c505",
   914 => x"78c148a6",
   915 => x"c548d0ff",
   916 => x"48d4ff78",
   917 => x"c478d5c1",
   918 => x"89c14966",
   919 => x"e4c131c6",
   920 => x"4abf97d8",
   921 => x"ffb07148",
   922 => x"ff7808d4",
   923 => x"78c448d0",
   924 => x"97f4e1c2",
   925 => x"99d049bf",
   926 => x"c587dd02",
   927 => x"48d4ff78",
   928 => x"c078d6c1",
   929 => x"48d4ff4a",
   930 => x"c178ffc3",
   931 => x"aae0c082",
   932 => x"ff87f204",
   933 => x"78c448d0",
   934 => x"c348d4ff",
   935 => x"d0ff78ff",
   936 => x"ff78c548",
   937 => x"d3c148d4",
   938 => x"ff78c178",
   939 => x"78c448d0",
   940 => x"06acb7c0",
   941 => x"c287cbc2",
   942 => x"4bbfc0e2",
   943 => x"737e748c",
   944 => x"ddc1029b",
   945 => x"4dc0c887",
   946 => x"abb7c08b",
   947 => x"c887c603",
   948 => x"c04da3c0",
   949 => x"f4e1c24b",
   950 => x"d049bf97",
   951 => x"87cf0299",
   952 => x"e1c21ec0",
   953 => x"dbeb49f8",
   954 => x"7086c487",
   955 => x"c287d84c",
   956 => x"c21ee4d4",
   957 => x"eb49f8e1",
   958 => x"4c7087ca",
   959 => x"d4c21e75",
   960 => x"f0fb49e4",
   961 => x"7486c887",
   962 => x"87c5059c",
   963 => x"cac148c0",
   964 => x"c21ec187",
   965 => x"e949f8e1",
   966 => x"86c487db",
   967 => x"fe059b73",
   968 => x"4c6e87e3",
   969 => x"06acb7c0",
   970 => x"e1c287d1",
   971 => x"78c048f8",
   972 => x"78c080d0",
   973 => x"e2c280f4",
   974 => x"c078bfc4",
   975 => x"fd01acb7",
   976 => x"d0ff87f5",
   977 => x"ff78c548",
   978 => x"d3c148d4",
   979 => x"ff78c078",
   980 => x"78c448d0",
   981 => x"c2c048c1",
   982 => x"f848c087",
   983 => x"264d268e",
   984 => x"264b264c",
   985 => x"5b5e0e4f",
   986 => x"fc0e5d5c",
   987 => x"c04d7186",
   988 => x"04ad4c4b",
   989 => x"c087e8c0",
   990 => x"741ed4f5",
   991 => x"87c4029c",
   992 => x"87c24ac0",
   993 => x"49724ac1",
   994 => x"c487feeb",
   995 => x"c17e7086",
   996 => x"c2056e83",
   997 => x"c14b7587",
   998 => x"06ab7584",
   999 => x"6e87d8ff",
  1000 => x"268efc48",
  1001 => x"264c264d",
  1002 => x"1e4f264b",
  1003 => x"66c44a71",
  1004 => x"7287c505",
  1005 => x"87e2f949",
  1006 => x"5e0e4f26",
  1007 => x"0e5d5c5b",
  1008 => x"4c7186fc",
  1009 => x"c291de49",
  1010 => x"714de4e2",
  1011 => x"026d9785",
  1012 => x"c287dcc1",
  1013 => x"49bfd4e2",
  1014 => x"fe718174",
  1015 => x"7e7087c7",
  1016 => x"c0029848",
  1017 => x"e2c287f2",
  1018 => x"4a704bd8",
  1019 => x"c4ff49cb",
  1020 => x"4b7487f1",
  1021 => x"e4c193cc",
  1022 => x"83c483e4",
  1023 => x"7bfcc0c1",
  1024 => x"c2c14974",
  1025 => x"7b7587d2",
  1026 => x"97dce4c1",
  1027 => x"c21e49bf",
  1028 => x"fe49d8e2",
  1029 => x"86c487d5",
  1030 => x"c1c14974",
  1031 => x"49c087fa",
  1032 => x"87d5c3c1",
  1033 => x"48f0e1c2",
  1034 => x"c04950c0",
  1035 => x"fc87c1e1",
  1036 => x"264d268e",
  1037 => x"264b264c",
  1038 => x"0000004f",
  1039 => x"64616f4c",
  1040 => x"2e676e69",
  1041 => x"00002e2e",
  1042 => x"61422080",
  1043 => x"00006b63",
  1044 => x"64616f4c",
  1045 => x"202e2a20",
  1046 => x"00000000",
  1047 => x"0000203a",
  1048 => x"61422080",
  1049 => x"00006b63",
  1050 => x"78452080",
  1051 => x"00007469",
  1052 => x"49204453",
  1053 => x"2e74696e",
  1054 => x"0000002e",
  1055 => x"00004b4f",
  1056 => x"544f4f42",
  1057 => x"20202020",
  1058 => x"004d4f52",
  1059 => x"711e731e",
  1060 => x"e2c2494b",
  1061 => x"7181bfd4",
  1062 => x"7087cafb",
  1063 => x"c4029a4a",
  1064 => x"dee54987",
  1065 => x"d4e2c287",
  1066 => x"7378c048",
  1067 => x"87fac149",
  1068 => x"4f264b26",
  1069 => x"711e731e",
  1070 => x"4aa3c44b",
  1071 => x"87d0c102",
  1072 => x"dc028ac1",
  1073 => x"c0028a87",
  1074 => x"058a87f2",
  1075 => x"c287d3c1",
  1076 => x"02bfd4e2",
  1077 => x"4887cbc1",
  1078 => x"e2c288c1",
  1079 => x"c1c158d8",
  1080 => x"d4e2c287",
  1081 => x"89c649bf",
  1082 => x"59d8e2c2",
  1083 => x"03a9b7c0",
  1084 => x"c287efc0",
  1085 => x"c048d4e2",
  1086 => x"87e6c078",
  1087 => x"bfd0e2c2",
  1088 => x"c287df02",
  1089 => x"48bfd4e2",
  1090 => x"e2c280c1",
  1091 => x"87d258d8",
  1092 => x"bfd0e2c2",
  1093 => x"c287cb02",
  1094 => x"48bfd4e2",
  1095 => x"e2c280c6",
  1096 => x"497358d8",
  1097 => x"4b2687c4",
  1098 => x"5e0e4f26",
  1099 => x"0e5d5c5b",
  1100 => x"a6d086f0",
  1101 => x"e4d4c259",
  1102 => x"c24cc04d",
  1103 => x"c148d0e2",
  1104 => x"48a6c878",
  1105 => x"7e7578c0",
  1106 => x"bfd4e2c2",
  1107 => x"06a8c048",
  1108 => x"c887c0c1",
  1109 => x"7e755ca6",
  1110 => x"48e4d4c2",
  1111 => x"f2c00298",
  1112 => x"4d66c487",
  1113 => x"1ed4f5c0",
  1114 => x"c40266cc",
  1115 => x"c24cc087",
  1116 => x"744cc187",
  1117 => x"87d1e449",
  1118 => x"7e7086c4",
  1119 => x"66c885c1",
  1120 => x"cc80c148",
  1121 => x"e2c258a6",
  1122 => x"03adbfd4",
  1123 => x"056e87c5",
  1124 => x"6e87d1ff",
  1125 => x"754cc04d",
  1126 => x"dcc3029d",
  1127 => x"d4f5c087",
  1128 => x"0266cc1e",
  1129 => x"a6c887c7",
  1130 => x"c578c048",
  1131 => x"48a6c887",
  1132 => x"66c878c1",
  1133 => x"87d1e349",
  1134 => x"7e7086c4",
  1135 => x"c2029848",
  1136 => x"cb4987e4",
  1137 => x"49699781",
  1138 => x"c10299d0",
  1139 => x"497487d4",
  1140 => x"e4c191cc",
  1141 => x"c2c181e4",
  1142 => x"81c879cc",
  1143 => x"7451ffc3",
  1144 => x"c291de49",
  1145 => x"714de4e2",
  1146 => x"97c1c285",
  1147 => x"49a5c17d",
  1148 => x"c251e0c0",
  1149 => x"bf97f4dc",
  1150 => x"c187d202",
  1151 => x"4ba5c284",
  1152 => x"4af4dcc2",
  1153 => x"fcfe49db",
  1154 => x"d9c187d9",
  1155 => x"49a5cd87",
  1156 => x"84c151c0",
  1157 => x"6e4ba5c2",
  1158 => x"fe49cb4a",
  1159 => x"c187c4fc",
  1160 => x"497487c4",
  1161 => x"e4c191cc",
  1162 => x"fec081e4",
  1163 => x"dcc279fa",
  1164 => x"02bf97f4",
  1165 => x"497487d8",
  1166 => x"84c191de",
  1167 => x"4be4e2c2",
  1168 => x"dcc28371",
  1169 => x"49dd4af4",
  1170 => x"87d7fbfe",
  1171 => x"4b7487d8",
  1172 => x"e2c293de",
  1173 => x"a3cb83e4",
  1174 => x"c151c049",
  1175 => x"4a6e7384",
  1176 => x"fafe49cb",
  1177 => x"66c887fd",
  1178 => x"cc80c148",
  1179 => x"acc758a6",
  1180 => x"87c5c003",
  1181 => x"e4fc056e",
  1182 => x"03acc787",
  1183 => x"c287e4c0",
  1184 => x"c048d0e2",
  1185 => x"cc497478",
  1186 => x"e4e4c191",
  1187 => x"fafec081",
  1188 => x"de497479",
  1189 => x"e4e2c291",
  1190 => x"c151c081",
  1191 => x"04acc784",
  1192 => x"c187dcff",
  1193 => x"c048c0e6",
  1194 => x"c180f750",
  1195 => x"c140d0cc",
  1196 => x"c878c8c1",
  1197 => x"f4c2c180",
  1198 => x"4966cc78",
  1199 => x"87d8f7c0",
  1200 => x"4d268ef0",
  1201 => x"4b264c26",
  1202 => x"731e4f26",
  1203 => x"494b711e",
  1204 => x"e4c191cc",
  1205 => x"a1c881e4",
  1206 => x"d8e4c14a",
  1207 => x"c9501248",
  1208 => x"f7c04aa1",
  1209 => x"501248f4",
  1210 => x"e4c181ca",
  1211 => x"501148dc",
  1212 => x"97dce4c1",
  1213 => x"c01e49bf",
  1214 => x"87eff249",
  1215 => x"e9f84973",
  1216 => x"268efc87",
  1217 => x"1e4f264b",
  1218 => x"f7c049c0",
  1219 => x"4f2687eb",
  1220 => x"494a711e",
  1221 => x"e4c191cc",
  1222 => x"81c881e4",
  1223 => x"48f0e1c2",
  1224 => x"f0c05011",
  1225 => x"f5fe49a2",
  1226 => x"49c087e2",
  1227 => x"2687c1d5",
  1228 => x"d4ff1e4f",
  1229 => x"7affc34a",
  1230 => x"c048d0ff",
  1231 => x"7ade78e1",
  1232 => x"c8487a71",
  1233 => x"7a7028b7",
  1234 => x"b7d04871",
  1235 => x"717a7028",
  1236 => x"28b7d848",
  1237 => x"d0ff7a70",
  1238 => x"78e0c048",
  1239 => x"5e0e4f26",
  1240 => x"0e5d5c5b",
  1241 => x"4d7186f4",
  1242 => x"c191cc49",
  1243 => x"c881e4e4",
  1244 => x"a1ca4aa1",
  1245 => x"48a6c47e",
  1246 => x"bfece1c2",
  1247 => x"bf976e78",
  1248 => x"4c66c44b",
  1249 => x"48122c73",
  1250 => x"7058a6cc",
  1251 => x"c984c19c",
  1252 => x"49699781",
  1253 => x"c204acb7",
  1254 => x"6e4cc087",
  1255 => x"c84abf97",
  1256 => x"31724966",
  1257 => x"66c4b9ff",
  1258 => x"72487499",
  1259 => x"b14a7030",
  1260 => x"59f0e1c2",
  1261 => x"87f9fd71",
  1262 => x"e2c21ec7",
  1263 => x"c11ebfcc",
  1264 => x"c21ee4e4",
  1265 => x"bf97f0e1",
  1266 => x"87f4c149",
  1267 => x"f3c04975",
  1268 => x"8ee887c6",
  1269 => x"4c264d26",
  1270 => x"4f264b26",
  1271 => x"711e731e",
  1272 => x"f9fd494b",
  1273 => x"fd497387",
  1274 => x"4b2687f4",
  1275 => x"731e4f26",
  1276 => x"c24b711e",
  1277 => x"d6024aa3",
  1278 => x"058ac187",
  1279 => x"c287e2c0",
  1280 => x"02bfcce2",
  1281 => x"c14887db",
  1282 => x"d0e2c288",
  1283 => x"c287d258",
  1284 => x"02bfd0e2",
  1285 => x"e2c287cb",
  1286 => x"c148bfcc",
  1287 => x"d0e2c280",
  1288 => x"c21ec758",
  1289 => x"1ebfcce2",
  1290 => x"1ee4e4c1",
  1291 => x"97f0e1c2",
  1292 => x"87cc49bf",
  1293 => x"f1c04973",
  1294 => x"8ef487de",
  1295 => x"4f264b26",
  1296 => x"5c5b5e0e",
  1297 => x"ccff0e5d",
  1298 => x"a6e8c086",
  1299 => x"48a6cc59",
  1300 => x"80c478c0",
  1301 => x"80c478c0",
  1302 => x"80c478c0",
  1303 => x"7866c8c1",
  1304 => x"78c180c4",
  1305 => x"78c180c4",
  1306 => x"48d0e2c2",
  1307 => x"dee078c1",
  1308 => x"87f8e087",
  1309 => x"7087cde0",
  1310 => x"adfbc04d",
  1311 => x"87f3c102",
  1312 => x"0566e4c0",
  1313 => x"c187e8c1",
  1314 => x"c44a66c4",
  1315 => x"c17e6a82",
  1316 => x"6e48d0c1",
  1317 => x"20412049",
  1318 => x"c1511041",
  1319 => x"c14866c4",
  1320 => x"6a78cacb",
  1321 => x"7581c749",
  1322 => x"66c4c151",
  1323 => x"c181c849",
  1324 => x"48a6dc51",
  1325 => x"c4c178c2",
  1326 => x"81c94966",
  1327 => x"c4c151c0",
  1328 => x"81ca4966",
  1329 => x"1ec151c0",
  1330 => x"496a1ed8",
  1331 => x"dfff81c8",
  1332 => x"86c887ee",
  1333 => x"4866c8c1",
  1334 => x"c701a8c0",
  1335 => x"48a6d487",
  1336 => x"87cf78c1",
  1337 => x"4866c8c1",
  1338 => x"a6dc88c1",
  1339 => x"ff87c458",
  1340 => x"7587f9de",
  1341 => x"f1cb029d",
  1342 => x"4866d487",
  1343 => x"a866ccc1",
  1344 => x"87e6cb03",
  1345 => x"ddff7ec0",
  1346 => x"4d7087fa",
  1347 => x"88c6c148",
  1348 => x"7058a6c8",
  1349 => x"d6c10298",
  1350 => x"88c94887",
  1351 => x"7058a6c8",
  1352 => x"d7c50298",
  1353 => x"88c14887",
  1354 => x"7058a6c8",
  1355 => x"f8c20298",
  1356 => x"88c34887",
  1357 => x"7058a6c8",
  1358 => x"87cf0298",
  1359 => x"c888c148",
  1360 => x"987058a6",
  1361 => x"87f4c402",
  1362 => x"c087fec9",
  1363 => x"dcff7ef0",
  1364 => x"4d7087f2",
  1365 => x"02adecc0",
  1366 => x"7e7587c2",
  1367 => x"02adecc0",
  1368 => x"dcff87cd",
  1369 => x"4d7087de",
  1370 => x"05adecc0",
  1371 => x"c087f3ff",
  1372 => x"c10566e4",
  1373 => x"ecc087ea",
  1374 => x"87c402ad",
  1375 => x"87c4dcff",
  1376 => x"1eca1ec0",
  1377 => x"cc4b66dc",
  1378 => x"66ccc193",
  1379 => x"4ca3c483",
  1380 => x"dcff496c",
  1381 => x"1ec187ea",
  1382 => x"496c1ede",
  1383 => x"87e0dcff",
  1384 => x"cbc186d0",
  1385 => x"a3c87bca",
  1386 => x"5166dc49",
  1387 => x"c049a3c9",
  1388 => x"ca5166e0",
  1389 => x"516e49a3",
  1390 => x"c14866dc",
  1391 => x"a6e0c080",
  1392 => x"4866d458",
  1393 => x"04a866d8",
  1394 => x"66d487cb",
  1395 => x"d880c148",
  1396 => x"fac758a6",
  1397 => x"4866d887",
  1398 => x"a6dc88c1",
  1399 => x"87efc758",
  1400 => x"87c8dbff",
  1401 => x"e6c74d70",
  1402 => x"fedcff87",
  1403 => x"58a6d087",
  1404 => x"06a866d0",
  1405 => x"a6d087c6",
  1406 => x"7866cc48",
  1407 => x"87ebdcff",
  1408 => x"05a8ecc0",
  1409 => x"c087f5c1",
  1410 => x"c10566e4",
  1411 => x"66d487e5",
  1412 => x"c191cc49",
  1413 => x"c48166c4",
  1414 => x"4c6a4aa1",
  1415 => x"cc4aa1c8",
  1416 => x"ccc15266",
  1417 => x"d9ff79d0",
  1418 => x"4d7087da",
  1419 => x"87da029d",
  1420 => x"02adfbc0",
  1421 => x"547587d4",
  1422 => x"87c8d9ff",
  1423 => x"029d4d70",
  1424 => x"c087c7c0",
  1425 => x"ff05adfb",
  1426 => x"e0c087ec",
  1427 => x"54c1c254",
  1428 => x"d47c97c0",
  1429 => x"66d84866",
  1430 => x"cbc004a8",
  1431 => x"4866d487",
  1432 => x"a6d880c1",
  1433 => x"87e7c558",
  1434 => x"c14866d8",
  1435 => x"58a6dc88",
  1436 => x"ff87dcc5",
  1437 => x"7087f5d8",
  1438 => x"87d3c54d",
  1439 => x"c04866cc",
  1440 => x"05a866e4",
  1441 => x"c087f4c4",
  1442 => x"c048a6e8",
  1443 => x"dadaff78",
  1444 => x"ff7e7087",
  1445 => x"c087d4da",
  1446 => x"c058a6f0",
  1447 => x"c005a8ec",
  1448 => x"48a687c7",
  1449 => x"c4c0786e",
  1450 => x"d7d7ff87",
  1451 => x"4966d487",
  1452 => x"c4c191cc",
  1453 => x"80714866",
  1454 => x"c458a6c8",
  1455 => x"82c84a66",
  1456 => x"ca4966c4",
  1457 => x"c0516e81",
  1458 => x"c14966ec",
  1459 => x"c1896e81",
  1460 => x"70307148",
  1461 => x"7189c149",
  1462 => x"e1c27a97",
  1463 => x"6e49bfec",
  1464 => x"4a6a9729",
  1465 => x"c0987148",
  1466 => x"c458a6f4",
  1467 => x"80c44866",
  1468 => x"c858a6cc",
  1469 => x"c04cbf66",
  1470 => x"cc4866e4",
  1471 => x"c002a866",
  1472 => x"7ec087c5",
  1473 => x"c187c2c0",
  1474 => x"c01e6e7e",
  1475 => x"49741ee0",
  1476 => x"87ecd6ff",
  1477 => x"4d7086c8",
  1478 => x"06adb7c0",
  1479 => x"7587d4c1",
  1480 => x"bf66c884",
  1481 => x"81e0c049",
  1482 => x"c14b8974",
  1483 => x"714adcc1",
  1484 => x"87efe7fe",
  1485 => x"7e7484c2",
  1486 => x"4866e8c0",
  1487 => x"ecc080c1",
  1488 => x"f0c058a6",
  1489 => x"81c14966",
  1490 => x"c002a970",
  1491 => x"4cc087c5",
  1492 => x"c187c2c0",
  1493 => x"cc1e744c",
  1494 => x"c049bf66",
  1495 => x"66c481e0",
  1496 => x"c81e7189",
  1497 => x"d5ff4966",
  1498 => x"86c887d6",
  1499 => x"01a8b7c0",
  1500 => x"c087c5ff",
  1501 => x"c00266e8",
  1502 => x"66c487d3",
  1503 => x"c081c949",
  1504 => x"c45166e8",
  1505 => x"cdc14866",
  1506 => x"cec078de",
  1507 => x"4966c487",
  1508 => x"51c281c9",
  1509 => x"c14866c4",
  1510 => x"d478dccf",
  1511 => x"66d84866",
  1512 => x"cbc004a8",
  1513 => x"4866d487",
  1514 => x"a6d880c1",
  1515 => x"87d1c058",
  1516 => x"c14866d8",
  1517 => x"58a6dc88",
  1518 => x"ff87c6c0",
  1519 => x"7087edd3",
  1520 => x"48a6cc4d",
  1521 => x"c6c078c0",
  1522 => x"dfd3ff87",
  1523 => x"c04d7087",
  1524 => x"c14866e0",
  1525 => x"a6e4c080",
  1526 => x"029d7558",
  1527 => x"d487cbc0",
  1528 => x"ccc14866",
  1529 => x"f404a866",
  1530 => x"66d487da",
  1531 => x"03a8c748",
  1532 => x"d487e1c0",
  1533 => x"e2c24c66",
  1534 => x"78c048d0",
  1535 => x"91cc4974",
  1536 => x"8166c4c1",
  1537 => x"6a4aa1c4",
  1538 => x"7952c04a",
  1539 => x"acc784c1",
  1540 => x"87e2ff04",
  1541 => x"0266e4c0",
  1542 => x"c187e2c0",
  1543 => x"c14966c4",
  1544 => x"c4c181d4",
  1545 => x"dcc14a66",
  1546 => x"c152c082",
  1547 => x"c179d0cc",
  1548 => x"c14966c4",
  1549 => x"c1c181d8",
  1550 => x"d6c079e0",
  1551 => x"66c4c187",
  1552 => x"81d4c149",
  1553 => x"4a66c4c1",
  1554 => x"c182d8c1",
  1555 => x"c17ae8c1",
  1556 => x"c179c7cc",
  1557 => x"c14966c4",
  1558 => x"cfc181e0",
  1559 => x"d1ff79ee",
  1560 => x"66d087c1",
  1561 => x"8eccff48",
  1562 => x"4c264d26",
  1563 => x"4f264b26",
  1564 => x"c21ec71e",
  1565 => x"1ebfcce2",
  1566 => x"1ee4e4c1",
  1567 => x"97f0e1c2",
  1568 => x"fbee49bf",
  1569 => x"e4e4c187",
  1570 => x"d9e1c049",
  1571 => x"268ef487",
  1572 => x"e4c11e4f",
  1573 => x"50c048d8",
  1574 => x"bfe0d3c2",
  1575 => x"f9d5ff49",
  1576 => x"2648c087",
  1577 => x"1e731e4f",
  1578 => x"c287c7c7",
  1579 => x"c048d8e2",
  1580 => x"48d4ff50",
  1581 => x"c178ffc3",
  1582 => x"fe49f0c1",
  1583 => x"fe87e8df",
  1584 => x"7087fdea",
  1585 => x"87cd0298",
  1586 => x"87f0f2fe",
  1587 => x"c4029870",
  1588 => x"c24ac187",
  1589 => x"724ac087",
  1590 => x"87c8029a",
  1591 => x"49fcc1c1",
  1592 => x"87c3dffe",
  1593 => x"48cce2c2",
  1594 => x"e1c278c0",
  1595 => x"50c048f0",
  1596 => x"87fcfd49",
  1597 => x"7087dafe",
  1598 => x"ce029b4b",
  1599 => x"c0e6c187",
  1600 => x"de49c75b",
  1601 => x"49c187d2",
  1602 => x"c287eedf",
  1603 => x"e1c087ed",
  1604 => x"87fa87cf",
  1605 => x"4f264b26",
  1606 => x"00000000",
  1607 => x"00000000",
  1608 => x"00000001",
  1609 => x"00000fba",
  1610 => x"000028a4",
  1611 => x"00000000",
  1612 => x"00000fba",
  1613 => x"000028c2",
  1614 => x"00000000",
  1615 => x"00000fba",
  1616 => x"000028e0",
  1617 => x"00000000",
  1618 => x"00000fba",
  1619 => x"000028fe",
  1620 => x"00000000",
  1621 => x"00000fba",
  1622 => x"0000291c",
  1623 => x"00000000",
  1624 => x"00000fba",
  1625 => x"0000293a",
  1626 => x"00000000",
  1627 => x"00000fba",
  1628 => x"00002958",
  1629 => x"00000000",
  1630 => x"00001310",
  1631 => x"00000000",
  1632 => x"00000000",
  1633 => x"000010b4",
  1634 => x"00000000",
  1635 => x"00000000",
  1636 => x"00001080",
  1637 => x"db86fc1e",
  1638 => x"fc7e7087",
  1639 => x"1e4f268e",
  1640 => x"c048f0fe",
  1641 => x"7909cd78",
  1642 => x"1e4f2609",
  1643 => x"49d4e6c1",
  1644 => x"4f2687ed",
  1645 => x"bff0fe1e",
  1646 => x"1e4f2648",
  1647 => x"c148f0fe",
  1648 => x"1e4f2678",
  1649 => x"c048f0fe",
  1650 => x"1e4f2678",
  1651 => x"52c04a71",
  1652 => x"0e4f2651",
  1653 => x"5d5c5b5e",
  1654 => x"7186f40e",
  1655 => x"7e6d974d",
  1656 => x"974ca5c1",
  1657 => x"a6c8486c",
  1658 => x"c4486e58",
  1659 => x"c505a866",
  1660 => x"c048ff87",
  1661 => x"caff87e6",
  1662 => x"49a5c287",
  1663 => x"714b6c97",
  1664 => x"6b974ba3",
  1665 => x"7e6c974b",
  1666 => x"80c1486e",
  1667 => x"c758a6c8",
  1668 => x"58a6cc98",
  1669 => x"fe7c9770",
  1670 => x"487387e1",
  1671 => x"4d268ef4",
  1672 => x"4b264c26",
  1673 => x"731e4f26",
  1674 => x"fe86f41e",
  1675 => x"bfe087d5",
  1676 => x"e0c0494b",
  1677 => x"c00299c0",
  1678 => x"4a7387ea",
  1679 => x"c29affc3",
  1680 => x"bf97cce6",
  1681 => x"cee6c249",
  1682 => x"c2517281",
  1683 => x"bf97cce6",
  1684 => x"c1486e7e",
  1685 => x"58a6c880",
  1686 => x"a6cc98c7",
  1687 => x"cce6c258",
  1688 => x"5066c848",
  1689 => x"7087cdfd",
  1690 => x"87cffd7e",
  1691 => x"4b268ef4",
  1692 => x"c21e4f26",
  1693 => x"fd49cce6",
  1694 => x"e8c187d1",
  1695 => x"defc49e6",
  1696 => x"87e8c487",
  1697 => x"5e0e4f26",
  1698 => x"0e5d5c5b",
  1699 => x"7e7186fc",
  1700 => x"c24dd4ff",
  1701 => x"fc49cce6",
  1702 => x"4b7087f9",
  1703 => x"04abb7c0",
  1704 => x"c387f5c2",
  1705 => x"c905abf0",
  1706 => x"e4edc187",
  1707 => x"c278c148",
  1708 => x"e0c387d6",
  1709 => x"87c905ab",
  1710 => x"48e8edc1",
  1711 => x"c7c278c1",
  1712 => x"e8edc187",
  1713 => x"87c602bf",
  1714 => x"4ca3c0c2",
  1715 => x"4c7387c2",
  1716 => x"bfe4edc1",
  1717 => x"87e0c002",
  1718 => x"b7c44974",
  1719 => x"edc19129",
  1720 => x"4a7481ec",
  1721 => x"92c29acf",
  1722 => x"307248c1",
  1723 => x"baff4a70",
  1724 => x"98694872",
  1725 => x"87db7970",
  1726 => x"b7c44974",
  1727 => x"edc19129",
  1728 => x"4a7481ec",
  1729 => x"92c29acf",
  1730 => x"307248c3",
  1731 => x"69484a70",
  1732 => x"6e7970b0",
  1733 => x"87e4c005",
  1734 => x"c848d0ff",
  1735 => x"7dc578e1",
  1736 => x"bfe8edc1",
  1737 => x"c387c302",
  1738 => x"edc17de0",
  1739 => x"c302bfe4",
  1740 => x"7df0c387",
  1741 => x"d0ff7d73",
  1742 => x"78e0c048",
  1743 => x"48e8edc1",
  1744 => x"edc178c0",
  1745 => x"78c048e4",
  1746 => x"49cce6c2",
  1747 => x"7087c4fa",
  1748 => x"abb7c04b",
  1749 => x"87cbfd03",
  1750 => x"8efc48c0",
  1751 => x"4c264d26",
  1752 => x"4f264b26",
  1753 => x"00000000",
  1754 => x"00000000",
  1755 => x"00000000",
  1756 => x"00000000",
  1757 => x"00000000",
  1758 => x"00000000",
  1759 => x"00000000",
  1760 => x"00000000",
  1761 => x"00000000",
  1762 => x"00000000",
  1763 => x"00000000",
  1764 => x"00000000",
  1765 => x"00000000",
  1766 => x"00000000",
  1767 => x"00000000",
  1768 => x"00000000",
  1769 => x"00000000",
  1770 => x"00000000",
  1771 => x"724ac01e",
  1772 => x"c191c449",
  1773 => x"c081eced",
  1774 => x"d082c179",
  1775 => x"ee04aab7",
  1776 => x"0e4f2687",
  1777 => x"5d5c5b5e",
  1778 => x"f74d710e",
  1779 => x"4a7587f5",
  1780 => x"922ab7c4",
  1781 => x"82ecedc1",
  1782 => x"9ccf4c75",
  1783 => x"496a94c2",
  1784 => x"c32b744b",
  1785 => x"7448c29b",
  1786 => x"ff4c7030",
  1787 => x"714874bc",
  1788 => x"f77a7098",
  1789 => x"487387c5",
  1790 => x"4c264d26",
  1791 => x"4f264b26",
  1792 => x"48d0ff1e",
  1793 => x"7178e1c8",
  1794 => x"08d4ff48",
  1795 => x"4866c478",
  1796 => x"7808d4ff",
  1797 => x"711e4f26",
  1798 => x"4966c44a",
  1799 => x"ff49721e",
  1800 => x"d0ff87de",
  1801 => x"78e0c048",
  1802 => x"4f268efc",
  1803 => x"711e731e",
  1804 => x"4966c84b",
  1805 => x"c14a731e",
  1806 => x"ff49a2e0",
  1807 => x"8efc87d8",
  1808 => x"4f264b26",
  1809 => x"48d0ff1e",
  1810 => x"7178c9c8",
  1811 => x"08d4ff48",
  1812 => x"1e4f2678",
  1813 => x"eb494a71",
  1814 => x"48d0ff87",
  1815 => x"4f2678c8",
  1816 => x"711e731e",
  1817 => x"e4e6c24b",
  1818 => x"87c302bf",
  1819 => x"ff87ebc2",
  1820 => x"c9c848d0",
  1821 => x"c0487378",
  1822 => x"d4ffb0e0",
  1823 => x"e6c27808",
  1824 => x"78c048d8",
  1825 => x"c50266c8",
  1826 => x"49ffc387",
  1827 => x"49c087c2",
  1828 => x"59e0e6c2",
  1829 => x"c60266cc",
  1830 => x"d5d5c587",
  1831 => x"cf87c44a",
  1832 => x"c24affff",
  1833 => x"c25ae4e6",
  1834 => x"c148e4e6",
  1835 => x"264b2678",
  1836 => x"5b5e0e4f",
  1837 => x"710e5d5c",
  1838 => x"e0e6c24d",
  1839 => x"9d754bbf",
  1840 => x"4987cb02",
  1841 => x"f1c191c8",
  1842 => x"82714ad8",
  1843 => x"f5c187c4",
  1844 => x"4cc04ad8",
  1845 => x"99734912",
  1846 => x"bfdce6c2",
  1847 => x"ffb87148",
  1848 => x"c17808d4",
  1849 => x"c8842bb7",
  1850 => x"e704acb7",
  1851 => x"d8e6c287",
  1852 => x"80c848bf",
  1853 => x"58dce6c2",
  1854 => x"4c264d26",
  1855 => x"4f264b26",
  1856 => x"711e731e",
  1857 => x"9a4a134b",
  1858 => x"7287cb02",
  1859 => x"87e1fe49",
  1860 => x"059a4a13",
  1861 => x"4b2687f5",
  1862 => x"c21e4f26",
  1863 => x"49bfd8e6",
  1864 => x"48d8e6c2",
  1865 => x"c478a1c1",
  1866 => x"03a9b7c0",
  1867 => x"d4ff87db",
  1868 => x"dce6c248",
  1869 => x"e6c278bf",
  1870 => x"c249bfd8",
  1871 => x"c148d8e6",
  1872 => x"c0c478a1",
  1873 => x"e504a9b7",
  1874 => x"48d0ff87",
  1875 => x"e6c278c8",
  1876 => x"78c048e4",
  1877 => x"00004f26",
  1878 => x"00000000",
  1879 => x"00000000",
  1880 => x"5f000000",
  1881 => x"0000005f",
  1882 => x"00030300",
  1883 => x"00000303",
  1884 => x"147f7f14",
  1885 => x"00147f7f",
  1886 => x"6b2e2400",
  1887 => x"00123a6b",
  1888 => x"18366a4c",
  1889 => x"0032566c",
  1890 => x"594f7e30",
  1891 => x"40683a77",
  1892 => x"07040000",
  1893 => x"00000003",
  1894 => x"3e1c0000",
  1895 => x"00004163",
  1896 => x"63410000",
  1897 => x"00001c3e",
  1898 => x"1c3e2a08",
  1899 => x"082a3e1c",
  1900 => x"3e080800",
  1901 => x"0008083e",
  1902 => x"e0800000",
  1903 => x"00000060",
  1904 => x"08080800",
  1905 => x"00080808",
  1906 => x"60000000",
  1907 => x"00000060",
  1908 => x"18306040",
  1909 => x"0103060c",
  1910 => x"597f3e00",
  1911 => x"003e7f4d",
  1912 => x"7f060400",
  1913 => x"0000007f",
  1914 => x"71634200",
  1915 => x"00464f59",
  1916 => x"49632200",
  1917 => x"00367f49",
  1918 => x"13161c18",
  1919 => x"00107f7f",
  1920 => x"45672700",
  1921 => x"00397d45",
  1922 => x"4b7e3c00",
  1923 => x"00307949",
  1924 => x"71010100",
  1925 => x"00070f79",
  1926 => x"497f3600",
  1927 => x"00367f49",
  1928 => x"494f0600",
  1929 => x"001e3f69",
  1930 => x"66000000",
  1931 => x"00000066",
  1932 => x"e6800000",
  1933 => x"00000066",
  1934 => x"14080800",
  1935 => x"00222214",
  1936 => x"14141400",
  1937 => x"00141414",
  1938 => x"14222200",
  1939 => x"00080814",
  1940 => x"51030200",
  1941 => x"00060f59",
  1942 => x"5d417f3e",
  1943 => x"001e1f55",
  1944 => x"097f7e00",
  1945 => x"007e7f09",
  1946 => x"497f7f00",
  1947 => x"00367f49",
  1948 => x"633e1c00",
  1949 => x"00414141",
  1950 => x"417f7f00",
  1951 => x"001c3e63",
  1952 => x"497f7f00",
  1953 => x"00414149",
  1954 => x"097f7f00",
  1955 => x"00010109",
  1956 => x"417f3e00",
  1957 => x"007a7b49",
  1958 => x"087f7f00",
  1959 => x"007f7f08",
  1960 => x"7f410000",
  1961 => x"0000417f",
  1962 => x"40602000",
  1963 => x"003f7f40",
  1964 => x"1c087f7f",
  1965 => x"00416336",
  1966 => x"407f7f00",
  1967 => x"00404040",
  1968 => x"0c067f7f",
  1969 => x"007f7f06",
  1970 => x"0c067f7f",
  1971 => x"007f7f18",
  1972 => x"417f3e00",
  1973 => x"003e7f41",
  1974 => x"097f7f00",
  1975 => x"00060f09",
  1976 => x"61417f3e",
  1977 => x"00407e7f",
  1978 => x"097f7f00",
  1979 => x"00667f19",
  1980 => x"4d6f2600",
  1981 => x"00327b59",
  1982 => x"7f010100",
  1983 => x"0001017f",
  1984 => x"407f3f00",
  1985 => x"003f7f40",
  1986 => x"703f0f00",
  1987 => x"000f3f70",
  1988 => x"18307f7f",
  1989 => x"007f7f30",
  1990 => x"1c366341",
  1991 => x"4163361c",
  1992 => x"7c060301",
  1993 => x"0103067c",
  1994 => x"4d597161",
  1995 => x"00414347",
  1996 => x"7f7f0000",
  1997 => x"00004141",
  1998 => x"0c060301",
  1999 => x"40603018",
  2000 => x"41410000",
  2001 => x"00007f7f",
  2002 => x"03060c08",
  2003 => x"00080c06",
  2004 => x"80808080",
  2005 => x"00808080",
  2006 => x"03000000",
  2007 => x"00000407",
  2008 => x"54742000",
  2009 => x"00787c54",
  2010 => x"447f7f00",
  2011 => x"00387c44",
  2012 => x"447c3800",
  2013 => x"00004444",
  2014 => x"447c3800",
  2015 => x"007f7f44",
  2016 => x"547c3800",
  2017 => x"00185c54",
  2018 => x"7f7e0400",
  2019 => x"00000505",
  2020 => x"a4bc1800",
  2021 => x"007cfca4",
  2022 => x"047f7f00",
  2023 => x"00787c04",
  2024 => x"3d000000",
  2025 => x"0000407d",
  2026 => x"80808000",
  2027 => x"00007dfd",
  2028 => x"107f7f00",
  2029 => x"00446c38",
  2030 => x"3f000000",
  2031 => x"0000407f",
  2032 => x"180c7c7c",
  2033 => x"00787c0c",
  2034 => x"047c7c00",
  2035 => x"00787c04",
  2036 => x"447c3800",
  2037 => x"00387c44",
  2038 => x"24fcfc00",
  2039 => x"00183c24",
  2040 => x"243c1800",
  2041 => x"00fcfc24",
  2042 => x"047c7c00",
  2043 => x"00080c04",
  2044 => x"545c4800",
  2045 => x"00207454",
  2046 => x"7f3f0400",
  2047 => x"00004444",
  2048 => x"407c3c00",
  2049 => x"007c7c40",
  2050 => x"603c1c00",
  2051 => x"001c3c60",
  2052 => x"30607c3c",
  2053 => x"003c7c60",
  2054 => x"10386c44",
  2055 => x"00446c38",
  2056 => x"e0bc1c00",
  2057 => x"001c3c60",
  2058 => x"74644400",
  2059 => x"00444c5c",
  2060 => x"3e080800",
  2061 => x"00414177",
  2062 => x"7f000000",
  2063 => x"0000007f",
  2064 => x"77414100",
  2065 => x"0008083e",
  2066 => x"03010102",
  2067 => x"00010202",
  2068 => x"7f7f7f7f",
  2069 => x"007f7f7f",
  2070 => x"1c1c0808",
  2071 => x"7f7f3e3e",
  2072 => x"3e3e7f7f",
  2073 => x"08081c1c",
  2074 => x"7c181000",
  2075 => x"0010187c",
  2076 => x"7c301000",
  2077 => x"0010307c",
  2078 => x"60603010",
  2079 => x"00061e78",
  2080 => x"183c6642",
  2081 => x"0042663c",
  2082 => x"c26a3878",
  2083 => x"00386cc6",
  2084 => x"60000060",
  2085 => x"00600000",
  2086 => x"5c5b5e0e",
  2087 => x"86fc0e5d",
  2088 => x"e6c27e71",
  2089 => x"c04cbfec",
  2090 => x"c41ec04b",
  2091 => x"c402ab66",
  2092 => x"c24dc087",
  2093 => x"754dc187",
  2094 => x"ee49731e",
  2095 => x"86c887e2",
  2096 => x"ef49e0c0",
  2097 => x"a4c487eb",
  2098 => x"f0496a4a",
  2099 => x"c9f187f2",
  2100 => x"c184cc87",
  2101 => x"abb7c883",
  2102 => x"87cdff04",
  2103 => x"4d268efc",
  2104 => x"4b264c26",
  2105 => x"711e4f26",
  2106 => x"f0e6c24a",
  2107 => x"f0e6c25a",
  2108 => x"4978c748",
  2109 => x"2687e1fe",
  2110 => x"1e731e4f",
  2111 => x"b7c04a71",
  2112 => x"87d303aa",
  2113 => x"bfe4d2c2",
  2114 => x"c187c405",
  2115 => x"c087c24b",
  2116 => x"e8d2c24b",
  2117 => x"c287c45b",
  2118 => x"fc5ae8d2",
  2119 => x"e4d2c248",
  2120 => x"c14a78bf",
  2121 => x"a2c0c19a",
  2122 => x"87e7ec49",
  2123 => x"4f264b26",
  2124 => x"c44a711e",
  2125 => x"49721e66",
  2126 => x"fc87f1eb",
  2127 => x"1e4f268e",
  2128 => x"c348d4ff",
  2129 => x"d0ff78ff",
  2130 => x"78e1c048",
  2131 => x"c148d4ff",
  2132 => x"c4487178",
  2133 => x"08d4ff30",
  2134 => x"48d0ff78",
  2135 => x"2678e0c0",
  2136 => x"5b5e0e4f",
  2137 => x"f00e5d5c",
  2138 => x"c87ec086",
  2139 => x"bfec48a6",
  2140 => x"c280fc78",
  2141 => x"78bfece6",
  2142 => x"bff4e6c2",
  2143 => x"4cbfe84d",
  2144 => x"bfe4d2c2",
  2145 => x"87fee349",
  2146 => x"f6e849c7",
  2147 => x"c2497087",
  2148 => x"87d00599",
  2149 => x"bfdcd2c2",
  2150 => x"c8b9ff49",
  2151 => x"99c19966",
  2152 => x"87c2c202",
  2153 => x"cb49e8cf",
  2154 => x"a6d087fe",
  2155 => x"e849c758",
  2156 => x"987087d1",
  2157 => x"c887c905",
  2158 => x"99c14966",
  2159 => x"87c6c102",
  2160 => x"c84b66cc",
  2161 => x"bfec48a6",
  2162 => x"e4d2c278",
  2163 => x"f5e249bf",
  2164 => x"cb497387",
  2165 => x"987087de",
  2166 => x"c287d702",
  2167 => x"49bfd8d2",
  2168 => x"d2c2b9c1",
  2169 => x"fd7159dc",
  2170 => x"e8cf87d5",
  2171 => x"87f8ca49",
  2172 => x"49c74b70",
  2173 => x"7087cce7",
  2174 => x"c6ff0598",
  2175 => x"4966c887",
  2176 => x"fe0599c1",
  2177 => x"d2c287fd",
  2178 => x"c14abfe4",
  2179 => x"e8d2c2ba",
  2180 => x"7a0afc5a",
  2181 => x"c19ac10a",
  2182 => x"e849a2c0",
  2183 => x"dac187f5",
  2184 => x"87dfe649",
  2185 => x"d2c27ec1",
  2186 => x"66c848dc",
  2187 => x"e4d2c278",
  2188 => x"c7c105bf",
  2189 => x"c0c0c887",
  2190 => x"d0d3c24b",
  2191 => x"49154d7e",
  2192 => x"87ffe549",
  2193 => x"c0029870",
  2194 => x"b47387c2",
  2195 => x"052bb7c1",
  2196 => x"7487ebff",
  2197 => x"99ffc349",
  2198 => x"49c01e71",
  2199 => x"7487d1fb",
  2200 => x"29b7c849",
  2201 => x"49c11e71",
  2202 => x"c887c5fb",
  2203 => x"49fdc386",
  2204 => x"c387d0e5",
  2205 => x"cae549fa",
  2206 => x"87fdc787",
  2207 => x"ffc34974",
  2208 => x"2cb7c899",
  2209 => x"9c74b471",
  2210 => x"87e5c002",
  2211 => x"ff48a6c8",
  2212 => x"c878bfc8",
  2213 => x"d2c24966",
  2214 => x"c289bfe0",
  2215 => x"c003a9e0",
  2216 => x"4cc087c5",
  2217 => x"c287d0c0",
  2218 => x"c848e0d2",
  2219 => x"c6c07866",
  2220 => x"e0d2c287",
  2221 => x"7478c048",
  2222 => x"0599c849",
  2223 => x"c387cec0",
  2224 => x"fee349f5",
  2225 => x"c2497087",
  2226 => x"e7c00299",
  2227 => x"f0e6c287",
  2228 => x"cac002bf",
  2229 => x"88c14887",
  2230 => x"58f4e6c2",
  2231 => x"c487d3c0",
  2232 => x"e0c14866",
  2233 => x"6e7e7080",
  2234 => x"c5c002bf",
  2235 => x"49ff4b87",
  2236 => x"7ec10f73",
  2237 => x"99c44974",
  2238 => x"87cec005",
  2239 => x"e349f2c3",
  2240 => x"497087c1",
  2241 => x"c00299c2",
  2242 => x"e6c287ed",
  2243 => x"487ebff0",
  2244 => x"03a8b7c7",
  2245 => x"6e87cbc0",
  2246 => x"c280c148",
  2247 => x"c058f4e6",
  2248 => x"66c487d3",
  2249 => x"80e0c148",
  2250 => x"bf6e7e70",
  2251 => x"87c5c002",
  2252 => x"7349fe4b",
  2253 => x"c37ec10f",
  2254 => x"c6e249fd",
  2255 => x"c2497087",
  2256 => x"e3c00299",
  2257 => x"f0e6c287",
  2258 => x"c9c002bf",
  2259 => x"f0e6c287",
  2260 => x"c078c048",
  2261 => x"66c487d0",
  2262 => x"82e0c14a",
  2263 => x"c5c0026a",
  2264 => x"49fd4b87",
  2265 => x"7ec10f73",
  2266 => x"e149fac3",
  2267 => x"497087d5",
  2268 => x"c00299c2",
  2269 => x"e6c287ea",
  2270 => x"c748bff0",
  2271 => x"c003a8b7",
  2272 => x"e6c287c9",
  2273 => x"78c748f0",
  2274 => x"c487d3c0",
  2275 => x"e0c14866",
  2276 => x"6e7e7080",
  2277 => x"c5c002bf",
  2278 => x"49fc4b87",
  2279 => x"7ec10f73",
  2280 => x"f0c34874",
  2281 => x"58a6cc98",
  2282 => x"c0059870",
  2283 => x"dac187ce",
  2284 => x"87cfe049",
  2285 => x"99c24970",
  2286 => x"87c1c202",
  2287 => x"c349e8cf",
  2288 => x"a6d087e6",
  2289 => x"e8e6c258",
  2290 => x"c250c048",
  2291 => x"bf97e8e6",
  2292 => x"87d9c105",
  2293 => x"c00566c8",
  2294 => x"dac187cd",
  2295 => x"e2dfff49",
  2296 => x"02987087",
  2297 => x"e887c6c1",
  2298 => x"c3494bbf",
  2299 => x"b7c899ff",
  2300 => x"c2b3712b",
  2301 => x"49bfe4d2",
  2302 => x"87cadaff",
  2303 => x"c24966cc",
  2304 => x"987087f2",
  2305 => x"87c6c002",
  2306 => x"48e8e6c2",
  2307 => x"e6c250c1",
  2308 => x"05bf97e8",
  2309 => x"7387d6c0",
  2310 => x"99f0c349",
  2311 => x"87c7ff05",
  2312 => x"ff49dac1",
  2313 => x"7087dcde",
  2314 => x"fafe0598",
  2315 => x"f0e6c287",
  2316 => x"cc4b49bf",
  2317 => x"8366c493",
  2318 => x"73714b6b",
  2319 => x"029d750f",
  2320 => x"6d87e9c0",
  2321 => x"87e4c002",
  2322 => x"ddff496d",
  2323 => x"497087f5",
  2324 => x"c00299c1",
  2325 => x"a5c487cb",
  2326 => x"f0e6c24b",
  2327 => x"4b6b49bf",
  2328 => x"0285c80f",
  2329 => x"6d87c5c0",
  2330 => x"87dcff05",
  2331 => x"c8c0026e",
  2332 => x"f0e6c287",
  2333 => x"dff049bf",
  2334 => x"268ef087",
  2335 => x"264c264d",
  2336 => x"004f264b",
  2337 => x"00000010",
  2338 => x"14111258",
  2339 => x"231c1b1d",
  2340 => x"9491595a",
  2341 => x"f4ebf2f5",
  2342 => x"00000000",
  2343 => x"00000000",
  2344 => x"00000000",
  2345 => x"00000000",
  2346 => x"ff4a711e",
  2347 => x"7249bfc8",
  2348 => x"4f2648a1",
  2349 => x"bfc8ff1e",
  2350 => x"c0c0fe89",
  2351 => x"a9c0c0c0",
  2352 => x"c087c401",
  2353 => x"c187c24a",
  2354 => x"2648724a",
  2355 => x"0000004f",
  2356 => x"11141258",
  2357 => x"231c1b1d",
  2358 => x"9194595a",
  2359 => x"f4ebf2f5",
  2360 => x"000024e4",
  2361 => x"4f545541",
  2362 => x"544f4f42",
  2363 => x"ab004247",
  2364 => x"ab000019",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
