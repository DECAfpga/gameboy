
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"f8",x"e6",x"c2",x"87"),
    12 => (x"48",x"c0",x"c8",x"4e"),
    13 => (x"d5",x"c1",x"28",x"c2"),
    14 => (x"ea",x"d6",x"e5",x"ea"),
    15 => (x"c1",x"46",x"71",x"49"),
    16 => (x"87",x"f9",x"01",x"88"),
    17 => (x"49",x"f8",x"e6",x"c2"),
    18 => (x"48",x"f4",x"d3",x"c2"),
    19 => (x"03",x"89",x"d0",x"89"),
    20 => (x"40",x"40",x"40",x"c0"),
    21 => (x"d0",x"87",x"f6",x"40"),
    22 => (x"50",x"c0",x"05",x"81"),
    23 => (x"f9",x"05",x"89",x"c1"),
    24 => (x"f3",x"d3",x"c2",x"87"),
    25 => (x"ef",x"d3",x"c2",x"4d"),
    26 => (x"02",x"ad",x"74",x"4c"),
    27 => (x"0f",x"24",x"87",x"c4"),
    28 => (x"e0",x"c1",x"87",x"f7"),
    29 => (x"d3",x"c2",x"87",x"ef"),
    30 => (x"d3",x"c2",x"4d",x"f3"),
    31 => (x"ad",x"74",x"4c",x"f3"),
    32 => (x"c4",x"87",x"c6",x"02"),
    33 => (x"f5",x"0f",x"6c",x"8c"),
    34 => (x"87",x"fd",x"00",x"87"),
    35 => (x"71",x"86",x"fc",x"1e"),
    36 => (x"49",x"c0",x"ff",x"4a"),
    37 => (x"c0",x"c4",x"48",x"69"),
    38 => (x"48",x"7e",x"70",x"98"),
    39 => (x"87",x"f4",x"02",x"98"),
    40 => (x"fc",x"48",x"79",x"72"),
    41 => (x"0e",x"4f",x"26",x"8e"),
    42 => (x"0e",x"5c",x"5b",x"5e"),
    43 => (x"4c",x"c0",x"4b",x"71"),
    44 => (x"02",x"9a",x"4a",x"13"),
    45 => (x"49",x"72",x"87",x"cd"),
    46 => (x"c1",x"87",x"d1",x"ff"),
    47 => (x"9a",x"4a",x"13",x"84"),
    48 => (x"74",x"87",x"f3",x"05"),
    49 => (x"26",x"4c",x"26",x"48"),
    50 => (x"1e",x"4f",x"26",x"4b"),
    51 => (x"1e",x"73",x"1e",x"72"),
    52 => (x"02",x"11",x"48",x"12"),
    53 => (x"c3",x"4b",x"87",x"ca"),
    54 => (x"73",x"9b",x"98",x"df"),
    55 => (x"87",x"f0",x"02",x"88"),
    56 => (x"4a",x"26",x"4b",x"26"),
    57 => (x"73",x"1e",x"4f",x"26"),
    58 => (x"c1",x"1e",x"72",x"1e"),
    59 => (x"87",x"ca",x"04",x"8b"),
    60 => (x"02",x"11",x"48",x"12"),
    61 => (x"02",x"88",x"87",x"c4"),
    62 => (x"4a",x"26",x"87",x"f1"),
    63 => (x"4f",x"26",x"4b",x"26"),
    64 => (x"73",x"1e",x"74",x"1e"),
    65 => (x"c1",x"1e",x"72",x"1e"),
    66 => (x"87",x"cf",x"04",x"8b"),
    67 => (x"02",x"11",x"48",x"12"),
    68 => (x"df",x"4c",x"87",x"c9"),
    69 => (x"88",x"74",x"9c",x"98"),
    70 => (x"26",x"87",x"ec",x"02"),
    71 => (x"26",x"4b",x"26",x"4a"),
    72 => (x"1e",x"4f",x"26",x"4c"),
    73 => (x"73",x"81",x"48",x"73"),
    74 => (x"87",x"c5",x"02",x"a9"),
    75 => (x"f6",x"05",x"53",x"12"),
    76 => (x"0e",x"4f",x"26",x"87"),
    77 => (x"0e",x"5c",x"5b",x"5e"),
    78 => (x"d4",x"ff",x"4a",x"71"),
    79 => (x"4b",x"66",x"cc",x"4c"),
    80 => (x"71",x"8b",x"c1",x"49"),
    81 => (x"87",x"ce",x"02",x"99"),
    82 => (x"6c",x"7c",x"ff",x"c3"),
    83 => (x"c1",x"49",x"73",x"52"),
    84 => (x"05",x"99",x"71",x"8b"),
    85 => (x"4c",x"26",x"87",x"f2"),
    86 => (x"4f",x"26",x"4b",x"26"),
    87 => (x"ff",x"1e",x"73",x"1e"),
    88 => (x"ff",x"c3",x"4b",x"d4"),
    89 => (x"c3",x"4a",x"6b",x"7b"),
    90 => (x"49",x"6b",x"7b",x"ff"),
    91 => (x"b1",x"72",x"32",x"c8"),
    92 => (x"6b",x"7b",x"ff",x"c3"),
    93 => (x"71",x"31",x"c8",x"4a"),
    94 => (x"7b",x"ff",x"c3",x"b2"),
    95 => (x"32",x"c8",x"49",x"6b"),
    96 => (x"48",x"71",x"b1",x"72"),
    97 => (x"4f",x"26",x"4b",x"26"),
    98 => (x"5c",x"5b",x"5e",x"0e"),
    99 => (x"4d",x"71",x"0e",x"5d"),
   100 => (x"75",x"4c",x"d4",x"ff"),
   101 => (x"98",x"ff",x"c3",x"48"),
   102 => (x"d3",x"c2",x"7c",x"70"),
   103 => (x"c8",x"05",x"bf",x"f4"),
   104 => (x"48",x"66",x"d0",x"87"),
   105 => (x"a6",x"d4",x"30",x"c9"),
   106 => (x"49",x"66",x"d0",x"58"),
   107 => (x"48",x"71",x"29",x"d8"),
   108 => (x"70",x"98",x"ff",x"c3"),
   109 => (x"49",x"66",x"d0",x"7c"),
   110 => (x"48",x"71",x"29",x"d0"),
   111 => (x"70",x"98",x"ff",x"c3"),
   112 => (x"49",x"66",x"d0",x"7c"),
   113 => (x"48",x"71",x"29",x"c8"),
   114 => (x"70",x"98",x"ff",x"c3"),
   115 => (x"48",x"66",x"d0",x"7c"),
   116 => (x"70",x"98",x"ff",x"c3"),
   117 => (x"d0",x"49",x"75",x"7c"),
   118 => (x"c3",x"48",x"71",x"29"),
   119 => (x"7c",x"70",x"98",x"ff"),
   120 => (x"f0",x"c9",x"4b",x"6c"),
   121 => (x"ff",x"c3",x"4a",x"ff"),
   122 => (x"87",x"cf",x"05",x"ab"),
   123 => (x"6c",x"7c",x"71",x"49"),
   124 => (x"02",x"8a",x"c1",x"4b"),
   125 => (x"ab",x"71",x"87",x"c5"),
   126 => (x"73",x"87",x"f2",x"02"),
   127 => (x"26",x"4d",x"26",x"48"),
   128 => (x"26",x"4b",x"26",x"4c"),
   129 => (x"49",x"c0",x"1e",x"4f"),
   130 => (x"c3",x"48",x"d4",x"ff"),
   131 => (x"81",x"c1",x"78",x"ff"),
   132 => (x"a9",x"b7",x"c8",x"c3"),
   133 => (x"26",x"87",x"f1",x"04"),
   134 => (x"5b",x"5e",x"0e",x"4f"),
   135 => (x"c0",x"0e",x"5d",x"5c"),
   136 => (x"f7",x"c1",x"f0",x"ff"),
   137 => (x"c0",x"c0",x"c1",x"4d"),
   138 => (x"4b",x"c0",x"c0",x"c0"),
   139 => (x"c4",x"87",x"d6",x"ff"),
   140 => (x"c0",x"4c",x"df",x"f8"),
   141 => (x"fd",x"49",x"75",x"1e"),
   142 => (x"86",x"c4",x"87",x"ce"),
   143 => (x"c0",x"05",x"a8",x"c1"),
   144 => (x"d4",x"ff",x"87",x"e5"),
   145 => (x"78",x"ff",x"c3",x"48"),
   146 => (x"e1",x"c0",x"1e",x"73"),
   147 => (x"49",x"e9",x"c1",x"f0"),
   148 => (x"c4",x"87",x"f5",x"fc"),
   149 => (x"05",x"98",x"70",x"86"),
   150 => (x"d4",x"ff",x"87",x"ca"),
   151 => (x"78",x"ff",x"c3",x"48"),
   152 => (x"87",x"cb",x"48",x"c1"),
   153 => (x"c1",x"87",x"de",x"fe"),
   154 => (x"c6",x"ff",x"05",x"8c"),
   155 => (x"26",x"48",x"c0",x"87"),
   156 => (x"26",x"4c",x"26",x"4d"),
   157 => (x"0e",x"4f",x"26",x"4b"),
   158 => (x"0e",x"5c",x"5b",x"5e"),
   159 => (x"c1",x"f0",x"ff",x"c0"),
   160 => (x"d4",x"ff",x"4c",x"c1"),
   161 => (x"78",x"ff",x"c3",x"48"),
   162 => (x"f8",x"49",x"fc",x"ca"),
   163 => (x"4b",x"d3",x"87",x"d9"),
   164 => (x"49",x"74",x"1e",x"c0"),
   165 => (x"c4",x"87",x"f1",x"fb"),
   166 => (x"05",x"98",x"70",x"86"),
   167 => (x"d4",x"ff",x"87",x"ca"),
   168 => (x"78",x"ff",x"c3",x"48"),
   169 => (x"87",x"cb",x"48",x"c1"),
   170 => (x"c1",x"87",x"da",x"fd"),
   171 => (x"df",x"ff",x"05",x"8b"),
   172 => (x"26",x"48",x"c0",x"87"),
   173 => (x"26",x"4b",x"26",x"4c"),
   174 => (x"00",x"00",x"00",x"4f"),
   175 => (x"00",x"44",x"4d",x"43"),
   176 => (x"43",x"48",x"44",x"53"),
   177 => (x"69",x"61",x"66",x"20"),
   178 => (x"00",x"0a",x"21",x"6c"),
   179 => (x"52",x"52",x"45",x"49"),
   180 => (x"00",x"00",x"00",x"00"),
   181 => (x"00",x"49",x"50",x"53"),
   182 => (x"74",x"69",x"72",x"57"),
   183 => (x"61",x"66",x"20",x"65"),
   184 => (x"64",x"65",x"6c",x"69"),
   185 => (x"5e",x"0e",x"00",x"0a"),
   186 => (x"0e",x"5d",x"5c",x"5b"),
   187 => (x"ff",x"4d",x"ff",x"c3"),
   188 => (x"d0",x"fc",x"4b",x"d4"),
   189 => (x"1e",x"ea",x"c6",x"87"),
   190 => (x"c1",x"f0",x"e1",x"c0"),
   191 => (x"c7",x"fa",x"49",x"c8"),
   192 => (x"c1",x"86",x"c4",x"87"),
   193 => (x"87",x"c8",x"02",x"a8"),
   194 => (x"c0",x"87",x"ec",x"fd"),
   195 => (x"87",x"e8",x"c1",x"48"),
   196 => (x"70",x"87",x"c9",x"f9"),
   197 => (x"ff",x"ff",x"cf",x"49"),
   198 => (x"a9",x"ea",x"c6",x"99"),
   199 => (x"fd",x"87",x"c8",x"02"),
   200 => (x"48",x"c0",x"87",x"d5"),
   201 => (x"75",x"87",x"d1",x"c1"),
   202 => (x"4c",x"f1",x"c0",x"7b"),
   203 => (x"70",x"87",x"ea",x"fb"),
   204 => (x"ec",x"c0",x"02",x"98"),
   205 => (x"c0",x"1e",x"c0",x"87"),
   206 => (x"fa",x"c1",x"f0",x"ff"),
   207 => (x"87",x"c8",x"f9",x"49"),
   208 => (x"98",x"70",x"86",x"c4"),
   209 => (x"75",x"87",x"da",x"05"),
   210 => (x"75",x"49",x"6b",x"7b"),
   211 => (x"75",x"7b",x"75",x"7b"),
   212 => (x"c1",x"7b",x"75",x"7b"),
   213 => (x"c4",x"02",x"99",x"c0"),
   214 => (x"db",x"48",x"c1",x"87"),
   215 => (x"d7",x"48",x"c0",x"87"),
   216 => (x"05",x"ac",x"c2",x"87"),
   217 => (x"c0",x"cb",x"87",x"ca"),
   218 => (x"87",x"fb",x"f4",x"49"),
   219 => (x"87",x"c8",x"48",x"c0"),
   220 => (x"fe",x"05",x"8c",x"c1"),
   221 => (x"48",x"c0",x"87",x"f6"),
   222 => (x"4c",x"26",x"4d",x"26"),
   223 => (x"4f",x"26",x"4b",x"26"),
   224 => (x"5c",x"5b",x"5e",x"0e"),
   225 => (x"d0",x"ff",x"0e",x"5d"),
   226 => (x"d0",x"e5",x"c0",x"4d"),
   227 => (x"c2",x"4c",x"c0",x"c1"),
   228 => (x"c1",x"48",x"f4",x"d3"),
   229 => (x"49",x"d4",x"cb",x"78"),
   230 => (x"c7",x"87",x"cc",x"f4"),
   231 => (x"f9",x"7d",x"c2",x"4b"),
   232 => (x"7d",x"c3",x"87",x"e3"),
   233 => (x"49",x"74",x"1e",x"c0"),
   234 => (x"c4",x"87",x"dd",x"f7"),
   235 => (x"05",x"a8",x"c1",x"86"),
   236 => (x"c2",x"4b",x"87",x"c1"),
   237 => (x"87",x"cb",x"05",x"ab"),
   238 => (x"f3",x"49",x"cc",x"cb"),
   239 => (x"48",x"c0",x"87",x"e9"),
   240 => (x"c1",x"87",x"f6",x"c0"),
   241 => (x"d4",x"ff",x"05",x"8b"),
   242 => (x"87",x"da",x"fc",x"87"),
   243 => (x"58",x"f8",x"d3",x"c2"),
   244 => (x"cd",x"05",x"98",x"70"),
   245 => (x"c0",x"1e",x"c1",x"87"),
   246 => (x"d0",x"c1",x"f0",x"ff"),
   247 => (x"87",x"e8",x"f6",x"49"),
   248 => (x"d4",x"ff",x"86",x"c4"),
   249 => (x"78",x"ff",x"c3",x"48"),
   250 => (x"c2",x"87",x"c3",x"c3"),
   251 => (x"c2",x"58",x"fc",x"d3"),
   252 => (x"48",x"d4",x"ff",x"7d"),
   253 => (x"c1",x"78",x"ff",x"c3"),
   254 => (x"26",x"4d",x"26",x"48"),
   255 => (x"26",x"4b",x"26",x"4c"),
   256 => (x"5b",x"5e",x"0e",x"4f"),
   257 => (x"fc",x"0e",x"5d",x"5c"),
   258 => (x"ff",x"4b",x"71",x"86"),
   259 => (x"7e",x"c0",x"4c",x"d4"),
   260 => (x"df",x"cd",x"ee",x"c5"),
   261 => (x"7c",x"ff",x"c3",x"4a"),
   262 => (x"fe",x"c3",x"48",x"6c"),
   263 => (x"f8",x"c0",x"05",x"a8"),
   264 => (x"73",x"4d",x"74",x"87"),
   265 => (x"87",x"cc",x"02",x"9b"),
   266 => (x"73",x"1e",x"66",x"d4"),
   267 => (x"87",x"c3",x"f4",x"49"),
   268 => (x"87",x"d4",x"86",x"c4"),
   269 => (x"c4",x"48",x"d0",x"ff"),
   270 => (x"66",x"d4",x"78",x"d1"),
   271 => (x"7d",x"ff",x"c3",x"4a"),
   272 => (x"f8",x"05",x"8a",x"c1"),
   273 => (x"5a",x"a6",x"d8",x"87"),
   274 => (x"7c",x"7c",x"ff",x"c3"),
   275 => (x"c5",x"05",x"9b",x"73"),
   276 => (x"48",x"d0",x"ff",x"87"),
   277 => (x"4a",x"c1",x"78",x"d0"),
   278 => (x"05",x"8a",x"c1",x"7e"),
   279 => (x"6e",x"87",x"f6",x"fe"),
   280 => (x"26",x"8e",x"fc",x"48"),
   281 => (x"26",x"4c",x"26",x"4d"),
   282 => (x"1e",x"4f",x"26",x"4b"),
   283 => (x"4a",x"71",x"1e",x"73"),
   284 => (x"d4",x"ff",x"4b",x"c0"),
   285 => (x"78",x"ff",x"c3",x"48"),
   286 => (x"c4",x"48",x"d0",x"ff"),
   287 => (x"d4",x"ff",x"78",x"c3"),
   288 => (x"78",x"ff",x"c3",x"48"),
   289 => (x"ff",x"c0",x"1e",x"72"),
   290 => (x"49",x"d1",x"c1",x"f0"),
   291 => (x"c4",x"87",x"f9",x"f3"),
   292 => (x"05",x"98",x"70",x"86"),
   293 => (x"c0",x"c8",x"87",x"d2"),
   294 => (x"49",x"66",x"cc",x"1e"),
   295 => (x"c4",x"87",x"e2",x"fd"),
   296 => (x"ff",x"4b",x"70",x"86"),
   297 => (x"78",x"c2",x"48",x"d0"),
   298 => (x"4b",x"26",x"48",x"73"),
   299 => (x"5e",x"0e",x"4f",x"26"),
   300 => (x"0e",x"5d",x"5c",x"5b"),
   301 => (x"ff",x"c0",x"1e",x"c0"),
   302 => (x"49",x"c9",x"c1",x"f0"),
   303 => (x"d2",x"87",x"c9",x"f3"),
   304 => (x"c4",x"d4",x"c2",x"1e"),
   305 => (x"87",x"f9",x"fc",x"49"),
   306 => (x"4c",x"c0",x"86",x"c8"),
   307 => (x"b7",x"d2",x"84",x"c1"),
   308 => (x"87",x"f8",x"04",x"ac"),
   309 => (x"97",x"c4",x"d4",x"c2"),
   310 => (x"c0",x"c3",x"49",x"bf"),
   311 => (x"a9",x"c0",x"c1",x"99"),
   312 => (x"87",x"e7",x"c0",x"05"),
   313 => (x"97",x"cb",x"d4",x"c2"),
   314 => (x"31",x"d0",x"49",x"bf"),
   315 => (x"97",x"cc",x"d4",x"c2"),
   316 => (x"32",x"c8",x"4a",x"bf"),
   317 => (x"d4",x"c2",x"b1",x"72"),
   318 => (x"4a",x"bf",x"97",x"cd"),
   319 => (x"cf",x"4c",x"71",x"b1"),
   320 => (x"9c",x"ff",x"ff",x"ff"),
   321 => (x"34",x"ca",x"84",x"c1"),
   322 => (x"c2",x"87",x"e7",x"c1"),
   323 => (x"bf",x"97",x"cd",x"d4"),
   324 => (x"c6",x"31",x"c1",x"49"),
   325 => (x"ce",x"d4",x"c2",x"99"),
   326 => (x"c7",x"4a",x"bf",x"97"),
   327 => (x"b1",x"72",x"2a",x"b7"),
   328 => (x"97",x"c9",x"d4",x"c2"),
   329 => (x"cf",x"4d",x"4a",x"bf"),
   330 => (x"ca",x"d4",x"c2",x"9d"),
   331 => (x"c3",x"4a",x"bf",x"97"),
   332 => (x"c2",x"32",x"ca",x"9a"),
   333 => (x"bf",x"97",x"cb",x"d4"),
   334 => (x"73",x"33",x"c2",x"4b"),
   335 => (x"cc",x"d4",x"c2",x"b2"),
   336 => (x"c3",x"4b",x"bf",x"97"),
   337 => (x"b7",x"c6",x"9b",x"c0"),
   338 => (x"c2",x"b2",x"73",x"2b"),
   339 => (x"71",x"48",x"c1",x"81"),
   340 => (x"c1",x"49",x"70",x"30"),
   341 => (x"70",x"30",x"75",x"48"),
   342 => (x"c1",x"4c",x"72",x"4d"),
   343 => (x"c8",x"94",x"71",x"84"),
   344 => (x"06",x"ad",x"b7",x"c0"),
   345 => (x"34",x"c1",x"87",x"cc"),
   346 => (x"c0",x"c8",x"2d",x"b7"),
   347 => (x"ff",x"01",x"ad",x"b7"),
   348 => (x"48",x"74",x"87",x"f4"),
   349 => (x"4c",x"26",x"4d",x"26"),
   350 => (x"4f",x"26",x"4b",x"26"),
   351 => (x"5c",x"5b",x"5e",x"0e"),
   352 => (x"86",x"fc",x"0e",x"5d"),
   353 => (x"48",x"ec",x"dc",x"c2"),
   354 => (x"d4",x"c2",x"78",x"c0"),
   355 => (x"49",x"c0",x"1e",x"e4"),
   356 => (x"c4",x"87",x"d8",x"fb"),
   357 => (x"05",x"98",x"70",x"86"),
   358 => (x"48",x"c0",x"87",x"c5"),
   359 => (x"c0",x"87",x"d1",x"c9"),
   360 => (x"e8",x"e1",x"c2",x"4d"),
   361 => (x"c2",x"78",x"c1",x"48"),
   362 => (x"c0",x"4a",x"da",x"d5"),
   363 => (x"c8",x"49",x"c8",x"e0"),
   364 => (x"87",x"f2",x"ec",x"4b"),
   365 => (x"c6",x"05",x"98",x"70"),
   366 => (x"e8",x"e1",x"c2",x"87"),
   367 => (x"c2",x"78",x"c0",x"48"),
   368 => (x"c0",x"4a",x"f6",x"d5"),
   369 => (x"c8",x"49",x"d4",x"e0"),
   370 => (x"87",x"da",x"ec",x"4b"),
   371 => (x"c6",x"05",x"98",x"70"),
   372 => (x"e8",x"e1",x"c2",x"87"),
   373 => (x"c2",x"78",x"c0",x"48"),
   374 => (x"02",x"bf",x"e8",x"e1"),
   375 => (x"c2",x"87",x"fd",x"c0"),
   376 => (x"4d",x"bf",x"ea",x"db"),
   377 => (x"9f",x"e2",x"dc",x"c2"),
   378 => (x"c5",x"48",x"7e",x"bf"),
   379 => (x"05",x"a8",x"ea",x"d6"),
   380 => (x"db",x"c2",x"87",x"c7"),
   381 => (x"ce",x"4d",x"bf",x"ea"),
   382 => (x"ca",x"48",x"6e",x"87"),
   383 => (x"02",x"a8",x"d5",x"e9"),
   384 => (x"48",x"c0",x"87",x"c5"),
   385 => (x"c2",x"87",x"e9",x"c7"),
   386 => (x"75",x"1e",x"e4",x"d4"),
   387 => (x"87",x"db",x"f9",x"49"),
   388 => (x"98",x"70",x"86",x"c4"),
   389 => (x"c0",x"87",x"c5",x"05"),
   390 => (x"87",x"d4",x"c7",x"48"),
   391 => (x"4a",x"f6",x"d5",x"c2"),
   392 => (x"49",x"e0",x"e0",x"c0"),
   393 => (x"fd",x"ea",x"4b",x"c8"),
   394 => (x"05",x"98",x"70",x"87"),
   395 => (x"dc",x"c2",x"87",x"c8"),
   396 => (x"78",x"c1",x"48",x"ec"),
   397 => (x"d5",x"c2",x"87",x"d8"),
   398 => (x"e0",x"c0",x"4a",x"da"),
   399 => (x"4b",x"c8",x"49",x"ec"),
   400 => (x"70",x"87",x"e3",x"ea"),
   401 => (x"c5",x"c0",x"02",x"98"),
   402 => (x"c6",x"48",x"c0",x"87"),
   403 => (x"dc",x"c2",x"87",x"e2"),
   404 => (x"49",x"bf",x"97",x"e2"),
   405 => (x"05",x"a9",x"d5",x"c1"),
   406 => (x"c2",x"87",x"cd",x"c0"),
   407 => (x"bf",x"97",x"e3",x"dc"),
   408 => (x"a9",x"ea",x"c2",x"49"),
   409 => (x"87",x"c5",x"c0",x"02"),
   410 => (x"c3",x"c6",x"48",x"c0"),
   411 => (x"e4",x"d4",x"c2",x"87"),
   412 => (x"48",x"7e",x"bf",x"97"),
   413 => (x"02",x"a8",x"e9",x"c3"),
   414 => (x"6e",x"87",x"ce",x"c0"),
   415 => (x"a8",x"eb",x"c3",x"48"),
   416 => (x"87",x"c5",x"c0",x"02"),
   417 => (x"e7",x"c5",x"48",x"c0"),
   418 => (x"ef",x"d4",x"c2",x"87"),
   419 => (x"99",x"49",x"bf",x"97"),
   420 => (x"87",x"cc",x"c0",x"05"),
   421 => (x"97",x"f0",x"d4",x"c2"),
   422 => (x"a9",x"c2",x"49",x"bf"),
   423 => (x"87",x"c5",x"c0",x"02"),
   424 => (x"cb",x"c5",x"48",x"c0"),
   425 => (x"f1",x"d4",x"c2",x"87"),
   426 => (x"c2",x"48",x"bf",x"97"),
   427 => (x"70",x"58",x"e8",x"dc"),
   428 => (x"88",x"c1",x"48",x"4c"),
   429 => (x"58",x"ec",x"dc",x"c2"),
   430 => (x"97",x"f2",x"d4",x"c2"),
   431 => (x"81",x"75",x"49",x"bf"),
   432 => (x"97",x"f3",x"d4",x"c2"),
   433 => (x"32",x"c8",x"4a",x"bf"),
   434 => (x"c2",x"7e",x"a1",x"72"),
   435 => (x"6e",x"48",x"c4",x"e1"),
   436 => (x"f4",x"d4",x"c2",x"78"),
   437 => (x"c2",x"48",x"bf",x"97"),
   438 => (x"c2",x"58",x"dc",x"e1"),
   439 => (x"02",x"bf",x"ec",x"dc"),
   440 => (x"c2",x"87",x"d2",x"c2"),
   441 => (x"df",x"4a",x"f6",x"d5"),
   442 => (x"4b",x"c8",x"49",x"fc"),
   443 => (x"70",x"87",x"f7",x"e7"),
   444 => (x"c5",x"c0",x"02",x"98"),
   445 => (x"c3",x"48",x"c0",x"87"),
   446 => (x"dc",x"c2",x"87",x"f6"),
   447 => (x"c2",x"4c",x"bf",x"e4"),
   448 => (x"c2",x"5c",x"d8",x"e1"),
   449 => (x"bf",x"97",x"c9",x"d5"),
   450 => (x"c2",x"31",x"c8",x"49"),
   451 => (x"bf",x"97",x"c8",x"d5"),
   452 => (x"c2",x"49",x"a1",x"4a"),
   453 => (x"bf",x"97",x"ca",x"d5"),
   454 => (x"72",x"32",x"d0",x"4a"),
   455 => (x"d5",x"c2",x"49",x"a1"),
   456 => (x"4a",x"bf",x"97",x"cb"),
   457 => (x"a1",x"72",x"32",x"d8"),
   458 => (x"e0",x"e1",x"c2",x"49"),
   459 => (x"d8",x"e1",x"c2",x"59"),
   460 => (x"e1",x"c2",x"91",x"bf"),
   461 => (x"c2",x"81",x"bf",x"c4"),
   462 => (x"c2",x"59",x"cc",x"e1"),
   463 => (x"bf",x"97",x"d1",x"d5"),
   464 => (x"c2",x"32",x"c8",x"4a"),
   465 => (x"bf",x"97",x"d0",x"d5"),
   466 => (x"c2",x"4a",x"a2",x"4b"),
   467 => (x"bf",x"97",x"d2",x"d5"),
   468 => (x"73",x"33",x"d0",x"4b"),
   469 => (x"d5",x"c2",x"4a",x"a2"),
   470 => (x"4b",x"bf",x"97",x"d3"),
   471 => (x"33",x"d8",x"9b",x"cf"),
   472 => (x"c2",x"4a",x"a2",x"73"),
   473 => (x"c2",x"5a",x"d0",x"e1"),
   474 => (x"c2",x"92",x"74",x"8a"),
   475 => (x"72",x"48",x"d0",x"e1"),
   476 => (x"c7",x"c1",x"78",x"a1"),
   477 => (x"f6",x"d4",x"c2",x"87"),
   478 => (x"c8",x"49",x"bf",x"97"),
   479 => (x"f5",x"d4",x"c2",x"31"),
   480 => (x"a1",x"4a",x"bf",x"97"),
   481 => (x"c7",x"31",x"c5",x"49"),
   482 => (x"29",x"c9",x"81",x"ff"),
   483 => (x"59",x"d8",x"e1",x"c2"),
   484 => (x"97",x"fb",x"d4",x"c2"),
   485 => (x"32",x"c8",x"4a",x"bf"),
   486 => (x"97",x"fa",x"d4",x"c2"),
   487 => (x"4a",x"a2",x"4b",x"bf"),
   488 => (x"5a",x"e0",x"e1",x"c2"),
   489 => (x"bf",x"d8",x"e1",x"c2"),
   490 => (x"c2",x"82",x"6e",x"92"),
   491 => (x"c2",x"5a",x"d4",x"e1"),
   492 => (x"c0",x"48",x"cc",x"e1"),
   493 => (x"c8",x"e1",x"c2",x"78"),
   494 => (x"78",x"a1",x"72",x"48"),
   495 => (x"48",x"e0",x"e1",x"c2"),
   496 => (x"bf",x"cc",x"e1",x"c2"),
   497 => (x"e4",x"e1",x"c2",x"78"),
   498 => (x"d0",x"e1",x"c2",x"48"),
   499 => (x"dc",x"c2",x"78",x"bf"),
   500 => (x"c0",x"02",x"bf",x"ec"),
   501 => (x"48",x"74",x"87",x"c9"),
   502 => (x"7e",x"70",x"30",x"c4"),
   503 => (x"c2",x"87",x"c9",x"c0"),
   504 => (x"48",x"bf",x"d4",x"e1"),
   505 => (x"7e",x"70",x"30",x"c4"),
   506 => (x"48",x"f0",x"dc",x"c2"),
   507 => (x"48",x"c1",x"78",x"6e"),
   508 => (x"4d",x"26",x"8e",x"fc"),
   509 => (x"4b",x"26",x"4c",x"26"),
   510 => (x"00",x"00",x"4f",x"26"),
   511 => (x"33",x"54",x"41",x"46"),
   512 => (x"20",x"20",x"20",x"32"),
   513 => (x"00",x"00",x"00",x"00"),
   514 => (x"31",x"54",x"41",x"46"),
   515 => (x"20",x"20",x"20",x"36"),
   516 => (x"00",x"00",x"00",x"00"),
   517 => (x"33",x"54",x"41",x"46"),
   518 => (x"20",x"20",x"20",x"32"),
   519 => (x"00",x"00",x"00",x"00"),
   520 => (x"33",x"54",x"41",x"46"),
   521 => (x"20",x"20",x"20",x"32"),
   522 => (x"00",x"00",x"00",x"00"),
   523 => (x"31",x"54",x"41",x"46"),
   524 => (x"20",x"20",x"20",x"36"),
   525 => (x"5b",x"5e",x"0e",x"00"),
   526 => (x"71",x"0e",x"5d",x"5c"),
   527 => (x"ec",x"dc",x"c2",x"4a"),
   528 => (x"87",x"cb",x"02",x"bf"),
   529 => (x"2b",x"c7",x"4b",x"72"),
   530 => (x"ff",x"c1",x"4d",x"72"),
   531 => (x"72",x"87",x"c9",x"9d"),
   532 => (x"72",x"2b",x"c8",x"4b"),
   533 => (x"9d",x"ff",x"c3",x"4d"),
   534 => (x"bf",x"c4",x"e1",x"c2"),
   535 => (x"c0",x"f2",x"c0",x"83"),
   536 => (x"d9",x"02",x"ab",x"bf"),
   537 => (x"c4",x"f2",x"c0",x"87"),
   538 => (x"e4",x"d4",x"c2",x"5b"),
   539 => (x"ef",x"49",x"73",x"1e"),
   540 => (x"86",x"c4",x"87",x"f9"),
   541 => (x"c5",x"05",x"98",x"70"),
   542 => (x"c0",x"48",x"c0",x"87"),
   543 => (x"dc",x"c2",x"87",x"e6"),
   544 => (x"d2",x"02",x"bf",x"ec"),
   545 => (x"c4",x"49",x"75",x"87"),
   546 => (x"e4",x"d4",x"c2",x"91"),
   547 => (x"cf",x"4c",x"69",x"81"),
   548 => (x"ff",x"ff",x"ff",x"ff"),
   549 => (x"75",x"87",x"cb",x"9c"),
   550 => (x"c2",x"91",x"c2",x"49"),
   551 => (x"9f",x"81",x"e4",x"d4"),
   552 => (x"48",x"74",x"4c",x"69"),
   553 => (x"4c",x"26",x"4d",x"26"),
   554 => (x"4f",x"26",x"4b",x"26"),
   555 => (x"5c",x"5b",x"5e",x"0e"),
   556 => (x"86",x"f4",x"0e",x"5d"),
   557 => (x"c8",x"59",x"a6",x"cc"),
   558 => (x"80",x"c8",x"48",x"66"),
   559 => (x"c0",x"48",x"7e",x"70"),
   560 => (x"49",x"c1",x"1e",x"78"),
   561 => (x"87",x"c1",x"c7",x"49"),
   562 => (x"4c",x"70",x"86",x"c4"),
   563 => (x"fb",x"c0",x"02",x"9c"),
   564 => (x"f4",x"dc",x"c2",x"87"),
   565 => (x"49",x"66",x"dc",x"4a"),
   566 => (x"87",x"ef",x"df",x"ff"),
   567 => (x"c0",x"02",x"98",x"70"),
   568 => (x"4a",x"74",x"87",x"ea"),
   569 => (x"cb",x"49",x"66",x"dc"),
   570 => (x"87",x"d4",x"e0",x"4b"),
   571 => (x"db",x"02",x"98",x"70"),
   572 => (x"74",x"1e",x"c0",x"87"),
   573 => (x"87",x"c4",x"02",x"9c"),
   574 => (x"87",x"c2",x"4d",x"c0"),
   575 => (x"49",x"75",x"4d",x"c1"),
   576 => (x"c4",x"87",x"c6",x"c6"),
   577 => (x"9c",x"4c",x"70",x"86"),
   578 => (x"87",x"c5",x"ff",x"05"),
   579 => (x"c1",x"02",x"9c",x"74"),
   580 => (x"a4",x"dc",x"87",x"d7"),
   581 => (x"69",x"48",x"6e",x"49"),
   582 => (x"49",x"a4",x"da",x"78"),
   583 => (x"c4",x"48",x"66",x"c8"),
   584 => (x"58",x"a6",x"c8",x"80"),
   585 => (x"c4",x"48",x"69",x"9f"),
   586 => (x"c2",x"78",x"08",x"66"),
   587 => (x"02",x"bf",x"ec",x"dc"),
   588 => (x"a4",x"d4",x"87",x"d2"),
   589 => (x"49",x"69",x"9f",x"49"),
   590 => (x"99",x"ff",x"ff",x"c0"),
   591 => (x"30",x"d0",x"48",x"71"),
   592 => (x"87",x"c2",x"7e",x"70"),
   593 => (x"48",x"6e",x"7e",x"c0"),
   594 => (x"80",x"bf",x"66",x"c4"),
   595 => (x"78",x"08",x"66",x"c4"),
   596 => (x"c0",x"48",x"66",x"c8"),
   597 => (x"49",x"66",x"c8",x"78"),
   598 => (x"66",x"c4",x"81",x"cc"),
   599 => (x"66",x"c8",x"79",x"bf"),
   600 => (x"c0",x"81",x"d0",x"49"),
   601 => (x"c2",x"48",x"c1",x"79"),
   602 => (x"f4",x"48",x"c0",x"87"),
   603 => (x"26",x"4d",x"26",x"8e"),
   604 => (x"26",x"4b",x"26",x"4c"),
   605 => (x"5b",x"5e",x"0e",x"4f"),
   606 => (x"71",x"0e",x"5d",x"5c"),
   607 => (x"4d",x"66",x"d0",x"4c"),
   608 => (x"72",x"49",x"6c",x"4a"),
   609 => (x"c2",x"b9",x"4d",x"a1"),
   610 => (x"4a",x"bf",x"e8",x"dc"),
   611 => (x"99",x"72",x"ba",x"ff"),
   612 => (x"c0",x"02",x"99",x"71"),
   613 => (x"a4",x"c4",x"87",x"e4"),
   614 => (x"fa",x"49",x"6b",x"4b"),
   615 => (x"7b",x"70",x"87",x"d7"),
   616 => (x"bf",x"e4",x"dc",x"c2"),
   617 => (x"71",x"81",x"6c",x"49"),
   618 => (x"c2",x"b9",x"75",x"7c"),
   619 => (x"4a",x"bf",x"e8",x"dc"),
   620 => (x"99",x"72",x"ba",x"ff"),
   621 => (x"ff",x"05",x"99",x"71"),
   622 => (x"7c",x"75",x"87",x"dc"),
   623 => (x"4c",x"26",x"4d",x"26"),
   624 => (x"4f",x"26",x"4b",x"26"),
   625 => (x"71",x"1e",x"73",x"1e"),
   626 => (x"c8",x"e1",x"c2",x"4b"),
   627 => (x"a3",x"c4",x"49",x"bf"),
   628 => (x"c2",x"4a",x"6a",x"4a"),
   629 => (x"e4",x"dc",x"c2",x"8a"),
   630 => (x"a1",x"72",x"92",x"bf"),
   631 => (x"e8",x"dc",x"c2",x"49"),
   632 => (x"9a",x"6b",x"4a",x"bf"),
   633 => (x"c0",x"49",x"a1",x"72"),
   634 => (x"c8",x"59",x"c4",x"f2"),
   635 => (x"e9",x"71",x"1e",x"66"),
   636 => (x"86",x"c4",x"87",x"f9"),
   637 => (x"c4",x"05",x"98",x"70"),
   638 => (x"c2",x"48",x"c0",x"87"),
   639 => (x"26",x"48",x"c1",x"87"),
   640 => (x"0e",x"4f",x"26",x"4b"),
   641 => (x"0e",x"5c",x"5b",x"5e"),
   642 => (x"4b",x"c0",x"4a",x"71"),
   643 => (x"c0",x"02",x"9a",x"72"),
   644 => (x"a2",x"da",x"87",x"e0"),
   645 => (x"4b",x"69",x"9f",x"49"),
   646 => (x"bf",x"ec",x"dc",x"c2"),
   647 => (x"d4",x"87",x"cf",x"02"),
   648 => (x"69",x"9f",x"49",x"a2"),
   649 => (x"ff",x"c0",x"4c",x"49"),
   650 => (x"34",x"d0",x"9c",x"ff"),
   651 => (x"4c",x"c0",x"87",x"c2"),
   652 => (x"9b",x"73",x"b3",x"74"),
   653 => (x"4a",x"87",x"df",x"02"),
   654 => (x"dc",x"c2",x"8a",x"c2"),
   655 => (x"92",x"49",x"bf",x"e4"),
   656 => (x"bf",x"c8",x"e1",x"c2"),
   657 => (x"c2",x"80",x"72",x"48"),
   658 => (x"71",x"58",x"e8",x"e1"),
   659 => (x"c2",x"30",x"c4",x"48"),
   660 => (x"c0",x"58",x"f4",x"dc"),
   661 => (x"e1",x"c2",x"87",x"e9"),
   662 => (x"c2",x"4b",x"bf",x"cc"),
   663 => (x"c2",x"48",x"e4",x"e1"),
   664 => (x"78",x"bf",x"d0",x"e1"),
   665 => (x"bf",x"ec",x"dc",x"c2"),
   666 => (x"c2",x"87",x"c9",x"02"),
   667 => (x"49",x"bf",x"e4",x"dc"),
   668 => (x"87",x"c7",x"31",x"c4"),
   669 => (x"bf",x"d4",x"e1",x"c2"),
   670 => (x"c2",x"31",x"c4",x"49"),
   671 => (x"c2",x"59",x"f4",x"dc"),
   672 => (x"26",x"5b",x"e4",x"e1"),
   673 => (x"26",x"4b",x"26",x"4c"),
   674 => (x"5b",x"5e",x"0e",x"4f"),
   675 => (x"f0",x"0e",x"5d",x"5c"),
   676 => (x"59",x"a6",x"c8",x"86"),
   677 => (x"ff",x"ff",x"ff",x"cf"),
   678 => (x"7e",x"c0",x"4c",x"f8"),
   679 => (x"d8",x"02",x"66",x"c4"),
   680 => (x"e0",x"d4",x"c2",x"87"),
   681 => (x"c2",x"78",x"c0",x"48"),
   682 => (x"c2",x"48",x"d8",x"d4"),
   683 => (x"78",x"bf",x"e4",x"e1"),
   684 => (x"48",x"dc",x"d4",x"c2"),
   685 => (x"bf",x"e0",x"e1",x"c2"),
   686 => (x"c1",x"dd",x"c2",x"78"),
   687 => (x"c2",x"50",x"c0",x"48"),
   688 => (x"49",x"bf",x"f0",x"dc"),
   689 => (x"bf",x"e0",x"d4",x"c2"),
   690 => (x"03",x"aa",x"71",x"4a"),
   691 => (x"72",x"87",x"cb",x"c4"),
   692 => (x"05",x"99",x"cf",x"49"),
   693 => (x"c0",x"87",x"e9",x"c0"),
   694 => (x"c2",x"48",x"c0",x"f2"),
   695 => (x"78",x"bf",x"d8",x"d4"),
   696 => (x"1e",x"e4",x"d4",x"c2"),
   697 => (x"bf",x"d8",x"d4",x"c2"),
   698 => (x"d8",x"d4",x"c2",x"49"),
   699 => (x"78",x"a1",x"c1",x"48"),
   700 => (x"87",x"f7",x"e5",x"71"),
   701 => (x"f1",x"c0",x"86",x"c4"),
   702 => (x"d4",x"c2",x"48",x"fc"),
   703 => (x"87",x"cc",x"78",x"e4"),
   704 => (x"bf",x"fc",x"f1",x"c0"),
   705 => (x"80",x"e0",x"c0",x"48"),
   706 => (x"58",x"c0",x"f2",x"c0"),
   707 => (x"bf",x"e0",x"d4",x"c2"),
   708 => (x"c2",x"80",x"c1",x"48"),
   709 => (x"27",x"58",x"e4",x"d4"),
   710 => (x"00",x"00",x"0c",x"7c"),
   711 => (x"4d",x"bf",x"97",x"bf"),
   712 => (x"e5",x"c2",x"02",x"9d"),
   713 => (x"ad",x"e5",x"c3",x"87"),
   714 => (x"87",x"de",x"c2",x"02"),
   715 => (x"bf",x"fc",x"f1",x"c0"),
   716 => (x"49",x"a3",x"cb",x"4b"),
   717 => (x"ac",x"cf",x"4c",x"11"),
   718 => (x"87",x"d2",x"c1",x"05"),
   719 => (x"99",x"df",x"49",x"75"),
   720 => (x"91",x"cd",x"89",x"c1"),
   721 => (x"81",x"f4",x"dc",x"c2"),
   722 => (x"12",x"4a",x"a3",x"c1"),
   723 => (x"4a",x"a3",x"c3",x"51"),
   724 => (x"a3",x"c5",x"51",x"12"),
   725 => (x"c7",x"51",x"12",x"4a"),
   726 => (x"51",x"12",x"4a",x"a3"),
   727 => (x"12",x"4a",x"a3",x"c9"),
   728 => (x"4a",x"a3",x"ce",x"51"),
   729 => (x"a3",x"d0",x"51",x"12"),
   730 => (x"d2",x"51",x"12",x"4a"),
   731 => (x"51",x"12",x"4a",x"a3"),
   732 => (x"12",x"4a",x"a3",x"d4"),
   733 => (x"4a",x"a3",x"d6",x"51"),
   734 => (x"a3",x"d8",x"51",x"12"),
   735 => (x"dc",x"51",x"12",x"4a"),
   736 => (x"51",x"12",x"4a",x"a3"),
   737 => (x"12",x"4a",x"a3",x"de"),
   738 => (x"c0",x"7e",x"c1",x"51"),
   739 => (x"49",x"74",x"87",x"fc"),
   740 => (x"c0",x"05",x"99",x"c8"),
   741 => (x"49",x"74",x"87",x"ed"),
   742 => (x"d3",x"05",x"99",x"d0"),
   743 => (x"66",x"e0",x"c0",x"87"),
   744 => (x"87",x"cc",x"c0",x"02"),
   745 => (x"e0",x"c0",x"49",x"73"),
   746 => (x"98",x"70",x"0f",x"66"),
   747 => (x"87",x"d3",x"c0",x"02"),
   748 => (x"c6",x"c0",x"05",x"6e"),
   749 => (x"f4",x"dc",x"c2",x"87"),
   750 => (x"c0",x"50",x"c0",x"48"),
   751 => (x"48",x"bf",x"fc",x"f1"),
   752 => (x"c2",x"87",x"e9",x"c2"),
   753 => (x"c0",x"48",x"c1",x"dd"),
   754 => (x"dc",x"c2",x"7e",x"50"),
   755 => (x"c2",x"49",x"bf",x"f0"),
   756 => (x"4a",x"bf",x"e0",x"d4"),
   757 => (x"fb",x"04",x"aa",x"71"),
   758 => (x"ff",x"cf",x"87",x"f5"),
   759 => (x"4c",x"f8",x"ff",x"ff"),
   760 => (x"bf",x"e4",x"e1",x"c2"),
   761 => (x"87",x"c8",x"c0",x"05"),
   762 => (x"bf",x"ec",x"dc",x"c2"),
   763 => (x"87",x"fa",x"c1",x"02"),
   764 => (x"bf",x"dc",x"d4",x"c2"),
   765 => (x"87",x"fd",x"f0",x"49"),
   766 => (x"58",x"e0",x"d4",x"c2"),
   767 => (x"c2",x"48",x"a6",x"c4"),
   768 => (x"78",x"bf",x"dc",x"d4"),
   769 => (x"bf",x"ec",x"dc",x"c2"),
   770 => (x"87",x"db",x"c0",x"02"),
   771 => (x"74",x"49",x"66",x"c4"),
   772 => (x"02",x"a9",x"74",x"99"),
   773 => (x"c8",x"87",x"c8",x"c0"),
   774 => (x"78",x"c0",x"48",x"a6"),
   775 => (x"c8",x"87",x"e7",x"c0"),
   776 => (x"78",x"c1",x"48",x"a6"),
   777 => (x"c4",x"87",x"df",x"c0"),
   778 => (x"ff",x"cf",x"49",x"66"),
   779 => (x"02",x"a9",x"99",x"f8"),
   780 => (x"cc",x"87",x"c8",x"c0"),
   781 => (x"78",x"c0",x"48",x"a6"),
   782 => (x"cc",x"87",x"c5",x"c0"),
   783 => (x"78",x"c1",x"48",x"a6"),
   784 => (x"cc",x"48",x"a6",x"c8"),
   785 => (x"66",x"c8",x"78",x"66"),
   786 => (x"87",x"de",x"c0",x"05"),
   787 => (x"c2",x"49",x"66",x"c4"),
   788 => (x"e4",x"dc",x"c2",x"89"),
   789 => (x"e1",x"c2",x"91",x"bf"),
   790 => (x"71",x"48",x"bf",x"c8"),
   791 => (x"dc",x"d4",x"c2",x"80"),
   792 => (x"e0",x"d4",x"c2",x"58"),
   793 => (x"f9",x"78",x"c0",x"48"),
   794 => (x"48",x"c0",x"87",x"d5"),
   795 => (x"ff",x"ff",x"ff",x"cf"),
   796 => (x"8e",x"f0",x"4c",x"f8"),
   797 => (x"4c",x"26",x"4d",x"26"),
   798 => (x"4f",x"26",x"4b",x"26"),
   799 => (x"00",x"00",x"00",x"00"),
   800 => (x"ff",x"ff",x"ff",x"ff"),
   801 => (x"48",x"d4",x"ff",x"1e"),
   802 => (x"68",x"78",x"ff",x"c3"),
   803 => (x"1e",x"4f",x"26",x"48"),
   804 => (x"c3",x"48",x"d4",x"ff"),
   805 => (x"d0",x"ff",x"78",x"ff"),
   806 => (x"78",x"e1",x"c0",x"48"),
   807 => (x"d4",x"48",x"d4",x"ff"),
   808 => (x"1e",x"4f",x"26",x"78"),
   809 => (x"c0",x"48",x"d0",x"ff"),
   810 => (x"4f",x"26",x"78",x"e0"),
   811 => (x"87",x"d4",x"ff",x"1e"),
   812 => (x"02",x"99",x"49",x"70"),
   813 => (x"fb",x"c0",x"87",x"c6"),
   814 => (x"87",x"f1",x"05",x"a9"),
   815 => (x"4f",x"26",x"48",x"71"),
   816 => (x"5c",x"5b",x"5e",x"0e"),
   817 => (x"c0",x"4b",x"71",x"0e"),
   818 => (x"87",x"f8",x"fe",x"4c"),
   819 => (x"02",x"99",x"49",x"70"),
   820 => (x"c0",x"87",x"f9",x"c0"),
   821 => (x"c0",x"02",x"a9",x"ec"),
   822 => (x"fb",x"c0",x"87",x"f2"),
   823 => (x"eb",x"c0",x"02",x"a9"),
   824 => (x"b7",x"66",x"cc",x"87"),
   825 => (x"87",x"c7",x"03",x"ac"),
   826 => (x"c2",x"02",x"66",x"d0"),
   827 => (x"71",x"53",x"71",x"87"),
   828 => (x"87",x"c2",x"02",x"99"),
   829 => (x"cb",x"fe",x"84",x"c1"),
   830 => (x"99",x"49",x"70",x"87"),
   831 => (x"c0",x"87",x"cd",x"02"),
   832 => (x"c7",x"02",x"a9",x"ec"),
   833 => (x"a9",x"fb",x"c0",x"87"),
   834 => (x"87",x"d5",x"ff",x"05"),
   835 => (x"c3",x"02",x"66",x"d0"),
   836 => (x"7b",x"97",x"c0",x"87"),
   837 => (x"05",x"a9",x"ec",x"c0"),
   838 => (x"4a",x"74",x"87",x"c4"),
   839 => (x"4a",x"74",x"87",x"c5"),
   840 => (x"72",x"8a",x"0a",x"c0"),
   841 => (x"26",x"4c",x"26",x"48"),
   842 => (x"1e",x"4f",x"26",x"4b"),
   843 => (x"70",x"87",x"d5",x"fd"),
   844 => (x"f0",x"c0",x"4a",x"49"),
   845 => (x"87",x"c9",x"04",x"aa"),
   846 => (x"01",x"aa",x"f9",x"c0"),
   847 => (x"f0",x"c0",x"87",x"c3"),
   848 => (x"aa",x"c1",x"c1",x"8a"),
   849 => (x"c1",x"87",x"c9",x"04"),
   850 => (x"c3",x"01",x"aa",x"da"),
   851 => (x"8a",x"f7",x"c0",x"87"),
   852 => (x"4f",x"26",x"48",x"72"),
   853 => (x"5c",x"5b",x"5e",x"0e"),
   854 => (x"86",x"f8",x"0e",x"5d"),
   855 => (x"7e",x"c0",x"4c",x"71"),
   856 => (x"c0",x"87",x"ec",x"fc"),
   857 => (x"f4",x"f7",x"c0",x"4b"),
   858 => (x"c0",x"49",x"bf",x"97"),
   859 => (x"87",x"cf",x"04",x"a9"),
   860 => (x"c1",x"87",x"f9",x"fc"),
   861 => (x"f4",x"f7",x"c0",x"83"),
   862 => (x"ab",x"49",x"bf",x"97"),
   863 => (x"c0",x"87",x"f1",x"06"),
   864 => (x"bf",x"97",x"f4",x"f7"),
   865 => (x"fb",x"87",x"cf",x"02"),
   866 => (x"49",x"70",x"87",x"fa"),
   867 => (x"87",x"c6",x"02",x"99"),
   868 => (x"05",x"a9",x"ec",x"c0"),
   869 => (x"4b",x"c0",x"87",x"f1"),
   870 => (x"70",x"87",x"e9",x"fb"),
   871 => (x"87",x"e4",x"fb",x"4d"),
   872 => (x"fb",x"58",x"a6",x"c8"),
   873 => (x"4a",x"70",x"87",x"de"),
   874 => (x"a4",x"c8",x"83",x"c1"),
   875 => (x"49",x"69",x"97",x"49"),
   876 => (x"87",x"da",x"05",x"ad"),
   877 => (x"97",x"49",x"a4",x"c9"),
   878 => (x"66",x"c4",x"49",x"69"),
   879 => (x"87",x"ce",x"05",x"a9"),
   880 => (x"97",x"49",x"a4",x"ca"),
   881 => (x"05",x"aa",x"49",x"69"),
   882 => (x"7e",x"c1",x"87",x"c4"),
   883 => (x"ec",x"c0",x"87",x"d0"),
   884 => (x"87",x"c6",x"02",x"ad"),
   885 => (x"05",x"ad",x"fb",x"c0"),
   886 => (x"4b",x"c0",x"87",x"c4"),
   887 => (x"02",x"6e",x"7e",x"c1"),
   888 => (x"fa",x"87",x"f5",x"fe"),
   889 => (x"48",x"73",x"87",x"fd"),
   890 => (x"4d",x"26",x"8e",x"f8"),
   891 => (x"4b",x"26",x"4c",x"26"),
   892 => (x"00",x"00",x"4f",x"26"),
   893 => (x"1e",x"73",x"1e",x"00"),
   894 => (x"c8",x"4b",x"d4",x"ff"),
   895 => (x"d0",x"ff",x"4a",x"66"),
   896 => (x"78",x"c5",x"c8",x"48"),
   897 => (x"c1",x"48",x"d4",x"ff"),
   898 => (x"7b",x"11",x"78",x"d4"),
   899 => (x"f9",x"05",x"8a",x"c1"),
   900 => (x"48",x"d0",x"ff",x"87"),
   901 => (x"4b",x"26",x"78",x"c4"),
   902 => (x"5e",x"0e",x"4f",x"26"),
   903 => (x"0e",x"5d",x"5c",x"5b"),
   904 => (x"7e",x"71",x"86",x"f8"),
   905 => (x"e1",x"c2",x"1e",x"6e"),
   906 => (x"ff",x"e9",x"49",x"f8"),
   907 => (x"70",x"86",x"c4",x"87"),
   908 => (x"e4",x"c4",x"02",x"98"),
   909 => (x"e0",x"e4",x"c1",x"87"),
   910 => (x"49",x"6e",x"4c",x"bf"),
   911 => (x"c8",x"87",x"d5",x"fc"),
   912 => (x"98",x"70",x"58",x"a6"),
   913 => (x"c4",x"87",x"c5",x"05"),
   914 => (x"78",x"c1",x"48",x"a6"),
   915 => (x"c5",x"48",x"d0",x"ff"),
   916 => (x"48",x"d4",x"ff",x"78"),
   917 => (x"c4",x"78",x"d5",x"c1"),
   918 => (x"89",x"c1",x"49",x"66"),
   919 => (x"e4",x"c1",x"31",x"c6"),
   920 => (x"4a",x"bf",x"97",x"d8"),
   921 => (x"ff",x"b0",x"71",x"48"),
   922 => (x"ff",x"78",x"08",x"d4"),
   923 => (x"78",x"c4",x"48",x"d0"),
   924 => (x"97",x"f4",x"e1",x"c2"),
   925 => (x"99",x"d0",x"49",x"bf"),
   926 => (x"c5",x"87",x"dd",x"02"),
   927 => (x"48",x"d4",x"ff",x"78"),
   928 => (x"c0",x"78",x"d6",x"c1"),
   929 => (x"48",x"d4",x"ff",x"4a"),
   930 => (x"c1",x"78",x"ff",x"c3"),
   931 => (x"aa",x"e0",x"c0",x"82"),
   932 => (x"ff",x"87",x"f2",x"04"),
   933 => (x"78",x"c4",x"48",x"d0"),
   934 => (x"c3",x"48",x"d4",x"ff"),
   935 => (x"d0",x"ff",x"78",x"ff"),
   936 => (x"ff",x"78",x"c5",x"48"),
   937 => (x"d3",x"c1",x"48",x"d4"),
   938 => (x"ff",x"78",x"c1",x"78"),
   939 => (x"78",x"c4",x"48",x"d0"),
   940 => (x"06",x"ac",x"b7",x"c0"),
   941 => (x"c2",x"87",x"cb",x"c2"),
   942 => (x"4b",x"bf",x"c0",x"e2"),
   943 => (x"73",x"7e",x"74",x"8c"),
   944 => (x"dd",x"c1",x"02",x"9b"),
   945 => (x"4d",x"c0",x"c8",x"87"),
   946 => (x"ab",x"b7",x"c0",x"8b"),
   947 => (x"c8",x"87",x"c6",x"03"),
   948 => (x"c0",x"4d",x"a3",x"c0"),
   949 => (x"f4",x"e1",x"c2",x"4b"),
   950 => (x"d0",x"49",x"bf",x"97"),
   951 => (x"87",x"cf",x"02",x"99"),
   952 => (x"e1",x"c2",x"1e",x"c0"),
   953 => (x"db",x"eb",x"49",x"f8"),
   954 => (x"70",x"86",x"c4",x"87"),
   955 => (x"c2",x"87",x"d8",x"4c"),
   956 => (x"c2",x"1e",x"e4",x"d4"),
   957 => (x"eb",x"49",x"f8",x"e1"),
   958 => (x"4c",x"70",x"87",x"ca"),
   959 => (x"d4",x"c2",x"1e",x"75"),
   960 => (x"f0",x"fb",x"49",x"e4"),
   961 => (x"74",x"86",x"c8",x"87"),
   962 => (x"87",x"c5",x"05",x"9c"),
   963 => (x"ca",x"c1",x"48",x"c0"),
   964 => (x"c2",x"1e",x"c1",x"87"),
   965 => (x"e9",x"49",x"f8",x"e1"),
   966 => (x"86",x"c4",x"87",x"db"),
   967 => (x"fe",x"05",x"9b",x"73"),
   968 => (x"4c",x"6e",x"87",x"e3"),
   969 => (x"06",x"ac",x"b7",x"c0"),
   970 => (x"e1",x"c2",x"87",x"d1"),
   971 => (x"78",x"c0",x"48",x"f8"),
   972 => (x"78",x"c0",x"80",x"d0"),
   973 => (x"e2",x"c2",x"80",x"f4"),
   974 => (x"c0",x"78",x"bf",x"c4"),
   975 => (x"fd",x"01",x"ac",x"b7"),
   976 => (x"d0",x"ff",x"87",x"f5"),
   977 => (x"ff",x"78",x"c5",x"48"),
   978 => (x"d3",x"c1",x"48",x"d4"),
   979 => (x"ff",x"78",x"c0",x"78"),
   980 => (x"78",x"c4",x"48",x"d0"),
   981 => (x"c2",x"c0",x"48",x"c1"),
   982 => (x"f8",x"48",x"c0",x"87"),
   983 => (x"26",x"4d",x"26",x"8e"),
   984 => (x"26",x"4b",x"26",x"4c"),
   985 => (x"5b",x"5e",x"0e",x"4f"),
   986 => (x"fc",x"0e",x"5d",x"5c"),
   987 => (x"c0",x"4d",x"71",x"86"),
   988 => (x"04",x"ad",x"4c",x"4b"),
   989 => (x"c0",x"87",x"e8",x"c0"),
   990 => (x"74",x"1e",x"d4",x"f5"),
   991 => (x"87",x"c4",x"02",x"9c"),
   992 => (x"87",x"c2",x"4a",x"c0"),
   993 => (x"49",x"72",x"4a",x"c1"),
   994 => (x"c4",x"87",x"fe",x"eb"),
   995 => (x"c1",x"7e",x"70",x"86"),
   996 => (x"c2",x"05",x"6e",x"83"),
   997 => (x"c1",x"4b",x"75",x"87"),
   998 => (x"06",x"ab",x"75",x"84"),
   999 => (x"6e",x"87",x"d8",x"ff"),
  1000 => (x"26",x"8e",x"fc",x"48"),
  1001 => (x"26",x"4c",x"26",x"4d"),
  1002 => (x"1e",x"4f",x"26",x"4b"),
  1003 => (x"66",x"c4",x"4a",x"71"),
  1004 => (x"72",x"87",x"c5",x"05"),
  1005 => (x"87",x"e2",x"f9",x"49"),
  1006 => (x"5e",x"0e",x"4f",x"26"),
  1007 => (x"0e",x"5d",x"5c",x"5b"),
  1008 => (x"4c",x"71",x"86",x"fc"),
  1009 => (x"c2",x"91",x"de",x"49"),
  1010 => (x"71",x"4d",x"e4",x"e2"),
  1011 => (x"02",x"6d",x"97",x"85"),
  1012 => (x"c2",x"87",x"dc",x"c1"),
  1013 => (x"49",x"bf",x"d4",x"e2"),
  1014 => (x"fe",x"71",x"81",x"74"),
  1015 => (x"7e",x"70",x"87",x"c7"),
  1016 => (x"c0",x"02",x"98",x"48"),
  1017 => (x"e2",x"c2",x"87",x"f2"),
  1018 => (x"4a",x"70",x"4b",x"d8"),
  1019 => (x"c4",x"ff",x"49",x"cb"),
  1020 => (x"4b",x"74",x"87",x"f1"),
  1021 => (x"e4",x"c1",x"93",x"cc"),
  1022 => (x"83",x"c4",x"83",x"e4"),
  1023 => (x"7b",x"fc",x"c0",x"c1"),
  1024 => (x"c2",x"c1",x"49",x"74"),
  1025 => (x"7b",x"75",x"87",x"d2"),
  1026 => (x"97",x"dc",x"e4",x"c1"),
  1027 => (x"c2",x"1e",x"49",x"bf"),
  1028 => (x"fe",x"49",x"d8",x"e2"),
  1029 => (x"86",x"c4",x"87",x"d5"),
  1030 => (x"c1",x"c1",x"49",x"74"),
  1031 => (x"49",x"c0",x"87",x"fa"),
  1032 => (x"87",x"d5",x"c3",x"c1"),
  1033 => (x"48",x"f0",x"e1",x"c2"),
  1034 => (x"c0",x"49",x"50",x"c0"),
  1035 => (x"fc",x"87",x"c1",x"e1"),
  1036 => (x"26",x"4d",x"26",x"8e"),
  1037 => (x"26",x"4b",x"26",x"4c"),
  1038 => (x"00",x"00",x"00",x"4f"),
  1039 => (x"64",x"61",x"6f",x"4c"),
  1040 => (x"2e",x"67",x"6e",x"69"),
  1041 => (x"00",x"00",x"2e",x"2e"),
  1042 => (x"61",x"42",x"20",x"80"),
  1043 => (x"00",x"00",x"6b",x"63"),
  1044 => (x"64",x"61",x"6f",x"4c"),
  1045 => (x"20",x"2e",x"2a",x"20"),
  1046 => (x"00",x"00",x"00",x"00"),
  1047 => (x"00",x"00",x"20",x"3a"),
  1048 => (x"61",x"42",x"20",x"80"),
  1049 => (x"00",x"00",x"6b",x"63"),
  1050 => (x"78",x"45",x"20",x"80"),
  1051 => (x"00",x"00",x"74",x"69"),
  1052 => (x"49",x"20",x"44",x"53"),
  1053 => (x"2e",x"74",x"69",x"6e"),
  1054 => (x"00",x"00",x"00",x"2e"),
  1055 => (x"00",x"00",x"4b",x"4f"),
  1056 => (x"54",x"4f",x"4f",x"42"),
  1057 => (x"20",x"20",x"20",x"20"),
  1058 => (x"00",x"4d",x"4f",x"52"),
  1059 => (x"71",x"1e",x"73",x"1e"),
  1060 => (x"e2",x"c2",x"49",x"4b"),
  1061 => (x"71",x"81",x"bf",x"d4"),
  1062 => (x"70",x"87",x"ca",x"fb"),
  1063 => (x"c4",x"02",x"9a",x"4a"),
  1064 => (x"de",x"e5",x"49",x"87"),
  1065 => (x"d4",x"e2",x"c2",x"87"),
  1066 => (x"73",x"78",x"c0",x"48"),
  1067 => (x"87",x"fa",x"c1",x"49"),
  1068 => (x"4f",x"26",x"4b",x"26"),
  1069 => (x"71",x"1e",x"73",x"1e"),
  1070 => (x"4a",x"a3",x"c4",x"4b"),
  1071 => (x"87",x"d0",x"c1",x"02"),
  1072 => (x"dc",x"02",x"8a",x"c1"),
  1073 => (x"c0",x"02",x"8a",x"87"),
  1074 => (x"05",x"8a",x"87",x"f2"),
  1075 => (x"c2",x"87",x"d3",x"c1"),
  1076 => (x"02",x"bf",x"d4",x"e2"),
  1077 => (x"48",x"87",x"cb",x"c1"),
  1078 => (x"e2",x"c2",x"88",x"c1"),
  1079 => (x"c1",x"c1",x"58",x"d8"),
  1080 => (x"d4",x"e2",x"c2",x"87"),
  1081 => (x"89",x"c6",x"49",x"bf"),
  1082 => (x"59",x"d8",x"e2",x"c2"),
  1083 => (x"03",x"a9",x"b7",x"c0"),
  1084 => (x"c2",x"87",x"ef",x"c0"),
  1085 => (x"c0",x"48",x"d4",x"e2"),
  1086 => (x"87",x"e6",x"c0",x"78"),
  1087 => (x"bf",x"d0",x"e2",x"c2"),
  1088 => (x"c2",x"87",x"df",x"02"),
  1089 => (x"48",x"bf",x"d4",x"e2"),
  1090 => (x"e2",x"c2",x"80",x"c1"),
  1091 => (x"87",x"d2",x"58",x"d8"),
  1092 => (x"bf",x"d0",x"e2",x"c2"),
  1093 => (x"c2",x"87",x"cb",x"02"),
  1094 => (x"48",x"bf",x"d4",x"e2"),
  1095 => (x"e2",x"c2",x"80",x"c6"),
  1096 => (x"49",x"73",x"58",x"d8"),
  1097 => (x"4b",x"26",x"87",x"c4"),
  1098 => (x"5e",x"0e",x"4f",x"26"),
  1099 => (x"0e",x"5d",x"5c",x"5b"),
  1100 => (x"a6",x"d0",x"86",x"f0"),
  1101 => (x"e4",x"d4",x"c2",x"59"),
  1102 => (x"c2",x"4c",x"c0",x"4d"),
  1103 => (x"c1",x"48",x"d0",x"e2"),
  1104 => (x"48",x"a6",x"c8",x"78"),
  1105 => (x"7e",x"75",x"78",x"c0"),
  1106 => (x"bf",x"d4",x"e2",x"c2"),
  1107 => (x"06",x"a8",x"c0",x"48"),
  1108 => (x"c8",x"87",x"c0",x"c1"),
  1109 => (x"7e",x"75",x"5c",x"a6"),
  1110 => (x"48",x"e4",x"d4",x"c2"),
  1111 => (x"f2",x"c0",x"02",x"98"),
  1112 => (x"4d",x"66",x"c4",x"87"),
  1113 => (x"1e",x"d4",x"f5",x"c0"),
  1114 => (x"c4",x"02",x"66",x"cc"),
  1115 => (x"c2",x"4c",x"c0",x"87"),
  1116 => (x"74",x"4c",x"c1",x"87"),
  1117 => (x"87",x"d1",x"e4",x"49"),
  1118 => (x"7e",x"70",x"86",x"c4"),
  1119 => (x"66",x"c8",x"85",x"c1"),
  1120 => (x"cc",x"80",x"c1",x"48"),
  1121 => (x"e2",x"c2",x"58",x"a6"),
  1122 => (x"03",x"ad",x"bf",x"d4"),
  1123 => (x"05",x"6e",x"87",x"c5"),
  1124 => (x"6e",x"87",x"d1",x"ff"),
  1125 => (x"75",x"4c",x"c0",x"4d"),
  1126 => (x"dc",x"c3",x"02",x"9d"),
  1127 => (x"d4",x"f5",x"c0",x"87"),
  1128 => (x"02",x"66",x"cc",x"1e"),
  1129 => (x"a6",x"c8",x"87",x"c7"),
  1130 => (x"c5",x"78",x"c0",x"48"),
  1131 => (x"48",x"a6",x"c8",x"87"),
  1132 => (x"66",x"c8",x"78",x"c1"),
  1133 => (x"87",x"d1",x"e3",x"49"),
  1134 => (x"7e",x"70",x"86",x"c4"),
  1135 => (x"c2",x"02",x"98",x"48"),
  1136 => (x"cb",x"49",x"87",x"e4"),
  1137 => (x"49",x"69",x"97",x"81"),
  1138 => (x"c1",x"02",x"99",x"d0"),
  1139 => (x"49",x"74",x"87",x"d4"),
  1140 => (x"e4",x"c1",x"91",x"cc"),
  1141 => (x"c2",x"c1",x"81",x"e4"),
  1142 => (x"81",x"c8",x"79",x"cc"),
  1143 => (x"74",x"51",x"ff",x"c3"),
  1144 => (x"c2",x"91",x"de",x"49"),
  1145 => (x"71",x"4d",x"e4",x"e2"),
  1146 => (x"97",x"c1",x"c2",x"85"),
  1147 => (x"49",x"a5",x"c1",x"7d"),
  1148 => (x"c2",x"51",x"e0",x"c0"),
  1149 => (x"bf",x"97",x"f4",x"dc"),
  1150 => (x"c1",x"87",x"d2",x"02"),
  1151 => (x"4b",x"a5",x"c2",x"84"),
  1152 => (x"4a",x"f4",x"dc",x"c2"),
  1153 => (x"fc",x"fe",x"49",x"db"),
  1154 => (x"d9",x"c1",x"87",x"d9"),
  1155 => (x"49",x"a5",x"cd",x"87"),
  1156 => (x"84",x"c1",x"51",x"c0"),
  1157 => (x"6e",x"4b",x"a5",x"c2"),
  1158 => (x"fe",x"49",x"cb",x"4a"),
  1159 => (x"c1",x"87",x"c4",x"fc"),
  1160 => (x"49",x"74",x"87",x"c4"),
  1161 => (x"e4",x"c1",x"91",x"cc"),
  1162 => (x"fe",x"c0",x"81",x"e4"),
  1163 => (x"dc",x"c2",x"79",x"fa"),
  1164 => (x"02",x"bf",x"97",x"f4"),
  1165 => (x"49",x"74",x"87",x"d8"),
  1166 => (x"84",x"c1",x"91",x"de"),
  1167 => (x"4b",x"e4",x"e2",x"c2"),
  1168 => (x"dc",x"c2",x"83",x"71"),
  1169 => (x"49",x"dd",x"4a",x"f4"),
  1170 => (x"87",x"d7",x"fb",x"fe"),
  1171 => (x"4b",x"74",x"87",x"d8"),
  1172 => (x"e2",x"c2",x"93",x"de"),
  1173 => (x"a3",x"cb",x"83",x"e4"),
  1174 => (x"c1",x"51",x"c0",x"49"),
  1175 => (x"4a",x"6e",x"73",x"84"),
  1176 => (x"fa",x"fe",x"49",x"cb"),
  1177 => (x"66",x"c8",x"87",x"fd"),
  1178 => (x"cc",x"80",x"c1",x"48"),
  1179 => (x"ac",x"c7",x"58",x"a6"),
  1180 => (x"87",x"c5",x"c0",x"03"),
  1181 => (x"e4",x"fc",x"05",x"6e"),
  1182 => (x"03",x"ac",x"c7",x"87"),
  1183 => (x"c2",x"87",x"e4",x"c0"),
  1184 => (x"c0",x"48",x"d0",x"e2"),
  1185 => (x"cc",x"49",x"74",x"78"),
  1186 => (x"e4",x"e4",x"c1",x"91"),
  1187 => (x"fa",x"fe",x"c0",x"81"),
  1188 => (x"de",x"49",x"74",x"79"),
  1189 => (x"e4",x"e2",x"c2",x"91"),
  1190 => (x"c1",x"51",x"c0",x"81"),
  1191 => (x"04",x"ac",x"c7",x"84"),
  1192 => (x"c1",x"87",x"dc",x"ff"),
  1193 => (x"c0",x"48",x"c0",x"e6"),
  1194 => (x"c1",x"80",x"f7",x"50"),
  1195 => (x"c1",x"40",x"d0",x"cc"),
  1196 => (x"c8",x"78",x"c8",x"c1"),
  1197 => (x"f4",x"c2",x"c1",x"80"),
  1198 => (x"49",x"66",x"cc",x"78"),
  1199 => (x"87",x"d8",x"f7",x"c0"),
  1200 => (x"4d",x"26",x"8e",x"f0"),
  1201 => (x"4b",x"26",x"4c",x"26"),
  1202 => (x"73",x"1e",x"4f",x"26"),
  1203 => (x"49",x"4b",x"71",x"1e"),
  1204 => (x"e4",x"c1",x"91",x"cc"),
  1205 => (x"a1",x"c8",x"81",x"e4"),
  1206 => (x"d8",x"e4",x"c1",x"4a"),
  1207 => (x"c9",x"50",x"12",x"48"),
  1208 => (x"f7",x"c0",x"4a",x"a1"),
  1209 => (x"50",x"12",x"48",x"f4"),
  1210 => (x"e4",x"c1",x"81",x"ca"),
  1211 => (x"50",x"11",x"48",x"dc"),
  1212 => (x"97",x"dc",x"e4",x"c1"),
  1213 => (x"c0",x"1e",x"49",x"bf"),
  1214 => (x"87",x"ef",x"f2",x"49"),
  1215 => (x"e9",x"f8",x"49",x"73"),
  1216 => (x"26",x"8e",x"fc",x"87"),
  1217 => (x"1e",x"4f",x"26",x"4b"),
  1218 => (x"f7",x"c0",x"49",x"c0"),
  1219 => (x"4f",x"26",x"87",x"eb"),
  1220 => (x"49",x"4a",x"71",x"1e"),
  1221 => (x"e4",x"c1",x"91",x"cc"),
  1222 => (x"81",x"c8",x"81",x"e4"),
  1223 => (x"48",x"f0",x"e1",x"c2"),
  1224 => (x"f0",x"c0",x"50",x"11"),
  1225 => (x"f5",x"fe",x"49",x"a2"),
  1226 => (x"49",x"c0",x"87",x"e2"),
  1227 => (x"26",x"87",x"c1",x"d5"),
  1228 => (x"d4",x"ff",x"1e",x"4f"),
  1229 => (x"7a",x"ff",x"c3",x"4a"),
  1230 => (x"c0",x"48",x"d0",x"ff"),
  1231 => (x"7a",x"de",x"78",x"e1"),
  1232 => (x"c8",x"48",x"7a",x"71"),
  1233 => (x"7a",x"70",x"28",x"b7"),
  1234 => (x"b7",x"d0",x"48",x"71"),
  1235 => (x"71",x"7a",x"70",x"28"),
  1236 => (x"28",x"b7",x"d8",x"48"),
  1237 => (x"d0",x"ff",x"7a",x"70"),
  1238 => (x"78",x"e0",x"c0",x"48"),
  1239 => (x"5e",x"0e",x"4f",x"26"),
  1240 => (x"0e",x"5d",x"5c",x"5b"),
  1241 => (x"4d",x"71",x"86",x"f4"),
  1242 => (x"c1",x"91",x"cc",x"49"),
  1243 => (x"c8",x"81",x"e4",x"e4"),
  1244 => (x"a1",x"ca",x"4a",x"a1"),
  1245 => (x"48",x"a6",x"c4",x"7e"),
  1246 => (x"bf",x"ec",x"e1",x"c2"),
  1247 => (x"bf",x"97",x"6e",x"78"),
  1248 => (x"4c",x"66",x"c4",x"4b"),
  1249 => (x"48",x"12",x"2c",x"73"),
  1250 => (x"70",x"58",x"a6",x"cc"),
  1251 => (x"c9",x"84",x"c1",x"9c"),
  1252 => (x"49",x"69",x"97",x"81"),
  1253 => (x"c2",x"04",x"ac",x"b7"),
  1254 => (x"6e",x"4c",x"c0",x"87"),
  1255 => (x"c8",x"4a",x"bf",x"97"),
  1256 => (x"31",x"72",x"49",x"66"),
  1257 => (x"66",x"c4",x"b9",x"ff"),
  1258 => (x"72",x"48",x"74",x"99"),
  1259 => (x"b1",x"4a",x"70",x"30"),
  1260 => (x"59",x"f0",x"e1",x"c2"),
  1261 => (x"87",x"f9",x"fd",x"71"),
  1262 => (x"e2",x"c2",x"1e",x"c7"),
  1263 => (x"c1",x"1e",x"bf",x"cc"),
  1264 => (x"c2",x"1e",x"e4",x"e4"),
  1265 => (x"bf",x"97",x"f0",x"e1"),
  1266 => (x"87",x"f4",x"c1",x"49"),
  1267 => (x"f3",x"c0",x"49",x"75"),
  1268 => (x"8e",x"e8",x"87",x"c6"),
  1269 => (x"4c",x"26",x"4d",x"26"),
  1270 => (x"4f",x"26",x"4b",x"26"),
  1271 => (x"71",x"1e",x"73",x"1e"),
  1272 => (x"f9",x"fd",x"49",x"4b"),
  1273 => (x"fd",x"49",x"73",x"87"),
  1274 => (x"4b",x"26",x"87",x"f4"),
  1275 => (x"73",x"1e",x"4f",x"26"),
  1276 => (x"c2",x"4b",x"71",x"1e"),
  1277 => (x"d6",x"02",x"4a",x"a3"),
  1278 => (x"05",x"8a",x"c1",x"87"),
  1279 => (x"c2",x"87",x"e2",x"c0"),
  1280 => (x"02",x"bf",x"cc",x"e2"),
  1281 => (x"c1",x"48",x"87",x"db"),
  1282 => (x"d0",x"e2",x"c2",x"88"),
  1283 => (x"c2",x"87",x"d2",x"58"),
  1284 => (x"02",x"bf",x"d0",x"e2"),
  1285 => (x"e2",x"c2",x"87",x"cb"),
  1286 => (x"c1",x"48",x"bf",x"cc"),
  1287 => (x"d0",x"e2",x"c2",x"80"),
  1288 => (x"c2",x"1e",x"c7",x"58"),
  1289 => (x"1e",x"bf",x"cc",x"e2"),
  1290 => (x"1e",x"e4",x"e4",x"c1"),
  1291 => (x"97",x"f0",x"e1",x"c2"),
  1292 => (x"87",x"cc",x"49",x"bf"),
  1293 => (x"f1",x"c0",x"49",x"73"),
  1294 => (x"8e",x"f4",x"87",x"de"),
  1295 => (x"4f",x"26",x"4b",x"26"),
  1296 => (x"5c",x"5b",x"5e",x"0e"),
  1297 => (x"cc",x"ff",x"0e",x"5d"),
  1298 => (x"a6",x"e8",x"c0",x"86"),
  1299 => (x"48",x"a6",x"cc",x"59"),
  1300 => (x"80",x"c4",x"78",x"c0"),
  1301 => (x"80",x"c4",x"78",x"c0"),
  1302 => (x"80",x"c4",x"78",x"c0"),
  1303 => (x"78",x"66",x"c8",x"c1"),
  1304 => (x"78",x"c1",x"80",x"c4"),
  1305 => (x"78",x"c1",x"80",x"c4"),
  1306 => (x"48",x"d0",x"e2",x"c2"),
  1307 => (x"de",x"e0",x"78",x"c1"),
  1308 => (x"87",x"f8",x"e0",x"87"),
  1309 => (x"70",x"87",x"cd",x"e0"),
  1310 => (x"ad",x"fb",x"c0",x"4d"),
  1311 => (x"87",x"f3",x"c1",x"02"),
  1312 => (x"05",x"66",x"e4",x"c0"),
  1313 => (x"c1",x"87",x"e8",x"c1"),
  1314 => (x"c4",x"4a",x"66",x"c4"),
  1315 => (x"c1",x"7e",x"6a",x"82"),
  1316 => (x"6e",x"48",x"d0",x"c1"),
  1317 => (x"20",x"41",x"20",x"49"),
  1318 => (x"c1",x"51",x"10",x"41"),
  1319 => (x"c1",x"48",x"66",x"c4"),
  1320 => (x"6a",x"78",x"ca",x"cb"),
  1321 => (x"75",x"81",x"c7",x"49"),
  1322 => (x"66",x"c4",x"c1",x"51"),
  1323 => (x"c1",x"81",x"c8",x"49"),
  1324 => (x"48",x"a6",x"dc",x"51"),
  1325 => (x"c4",x"c1",x"78",x"c2"),
  1326 => (x"81",x"c9",x"49",x"66"),
  1327 => (x"c4",x"c1",x"51",x"c0"),
  1328 => (x"81",x"ca",x"49",x"66"),
  1329 => (x"1e",x"c1",x"51",x"c0"),
  1330 => (x"49",x"6a",x"1e",x"d8"),
  1331 => (x"df",x"ff",x"81",x"c8"),
  1332 => (x"86",x"c8",x"87",x"ee"),
  1333 => (x"48",x"66",x"c8",x"c1"),
  1334 => (x"c7",x"01",x"a8",x"c0"),
  1335 => (x"48",x"a6",x"d4",x"87"),
  1336 => (x"87",x"cf",x"78",x"c1"),
  1337 => (x"48",x"66",x"c8",x"c1"),
  1338 => (x"a6",x"dc",x"88",x"c1"),
  1339 => (x"ff",x"87",x"c4",x"58"),
  1340 => (x"75",x"87",x"f9",x"de"),
  1341 => (x"f1",x"cb",x"02",x"9d"),
  1342 => (x"48",x"66",x"d4",x"87"),
  1343 => (x"a8",x"66",x"cc",x"c1"),
  1344 => (x"87",x"e6",x"cb",x"03"),
  1345 => (x"dd",x"ff",x"7e",x"c0"),
  1346 => (x"4d",x"70",x"87",x"fa"),
  1347 => (x"88",x"c6",x"c1",x"48"),
  1348 => (x"70",x"58",x"a6",x"c8"),
  1349 => (x"d6",x"c1",x"02",x"98"),
  1350 => (x"88",x"c9",x"48",x"87"),
  1351 => (x"70",x"58",x"a6",x"c8"),
  1352 => (x"d7",x"c5",x"02",x"98"),
  1353 => (x"88",x"c1",x"48",x"87"),
  1354 => (x"70",x"58",x"a6",x"c8"),
  1355 => (x"f8",x"c2",x"02",x"98"),
  1356 => (x"88",x"c3",x"48",x"87"),
  1357 => (x"70",x"58",x"a6",x"c8"),
  1358 => (x"87",x"cf",x"02",x"98"),
  1359 => (x"c8",x"88",x"c1",x"48"),
  1360 => (x"98",x"70",x"58",x"a6"),
  1361 => (x"87",x"f4",x"c4",x"02"),
  1362 => (x"c0",x"87",x"fe",x"c9"),
  1363 => (x"dc",x"ff",x"7e",x"f0"),
  1364 => (x"4d",x"70",x"87",x"f2"),
  1365 => (x"02",x"ad",x"ec",x"c0"),
  1366 => (x"7e",x"75",x"87",x"c2"),
  1367 => (x"02",x"ad",x"ec",x"c0"),
  1368 => (x"dc",x"ff",x"87",x"cd"),
  1369 => (x"4d",x"70",x"87",x"de"),
  1370 => (x"05",x"ad",x"ec",x"c0"),
  1371 => (x"c0",x"87",x"f3",x"ff"),
  1372 => (x"c1",x"05",x"66",x"e4"),
  1373 => (x"ec",x"c0",x"87",x"ea"),
  1374 => (x"87",x"c4",x"02",x"ad"),
  1375 => (x"87",x"c4",x"dc",x"ff"),
  1376 => (x"1e",x"ca",x"1e",x"c0"),
  1377 => (x"cc",x"4b",x"66",x"dc"),
  1378 => (x"66",x"cc",x"c1",x"93"),
  1379 => (x"4c",x"a3",x"c4",x"83"),
  1380 => (x"dc",x"ff",x"49",x"6c"),
  1381 => (x"1e",x"c1",x"87",x"ea"),
  1382 => (x"49",x"6c",x"1e",x"de"),
  1383 => (x"87",x"e0",x"dc",x"ff"),
  1384 => (x"cb",x"c1",x"86",x"d0"),
  1385 => (x"a3",x"c8",x"7b",x"ca"),
  1386 => (x"51",x"66",x"dc",x"49"),
  1387 => (x"c0",x"49",x"a3",x"c9"),
  1388 => (x"ca",x"51",x"66",x"e0"),
  1389 => (x"51",x"6e",x"49",x"a3"),
  1390 => (x"c1",x"48",x"66",x"dc"),
  1391 => (x"a6",x"e0",x"c0",x"80"),
  1392 => (x"48",x"66",x"d4",x"58"),
  1393 => (x"04",x"a8",x"66",x"d8"),
  1394 => (x"66",x"d4",x"87",x"cb"),
  1395 => (x"d8",x"80",x"c1",x"48"),
  1396 => (x"fa",x"c7",x"58",x"a6"),
  1397 => (x"48",x"66",x"d8",x"87"),
  1398 => (x"a6",x"dc",x"88",x"c1"),
  1399 => (x"87",x"ef",x"c7",x"58"),
  1400 => (x"87",x"c8",x"db",x"ff"),
  1401 => (x"e6",x"c7",x"4d",x"70"),
  1402 => (x"fe",x"dc",x"ff",x"87"),
  1403 => (x"58",x"a6",x"d0",x"87"),
  1404 => (x"06",x"a8",x"66",x"d0"),
  1405 => (x"a6",x"d0",x"87",x"c6"),
  1406 => (x"78",x"66",x"cc",x"48"),
  1407 => (x"87",x"eb",x"dc",x"ff"),
  1408 => (x"05",x"a8",x"ec",x"c0"),
  1409 => (x"c0",x"87",x"f5",x"c1"),
  1410 => (x"c1",x"05",x"66",x"e4"),
  1411 => (x"66",x"d4",x"87",x"e5"),
  1412 => (x"c1",x"91",x"cc",x"49"),
  1413 => (x"c4",x"81",x"66",x"c4"),
  1414 => (x"4c",x"6a",x"4a",x"a1"),
  1415 => (x"cc",x"4a",x"a1",x"c8"),
  1416 => (x"cc",x"c1",x"52",x"66"),
  1417 => (x"d9",x"ff",x"79",x"d0"),
  1418 => (x"4d",x"70",x"87",x"da"),
  1419 => (x"87",x"da",x"02",x"9d"),
  1420 => (x"02",x"ad",x"fb",x"c0"),
  1421 => (x"54",x"75",x"87",x"d4"),
  1422 => (x"87",x"c8",x"d9",x"ff"),
  1423 => (x"02",x"9d",x"4d",x"70"),
  1424 => (x"c0",x"87",x"c7",x"c0"),
  1425 => (x"ff",x"05",x"ad",x"fb"),
  1426 => (x"e0",x"c0",x"87",x"ec"),
  1427 => (x"54",x"c1",x"c2",x"54"),
  1428 => (x"d4",x"7c",x"97",x"c0"),
  1429 => (x"66",x"d8",x"48",x"66"),
  1430 => (x"cb",x"c0",x"04",x"a8"),
  1431 => (x"48",x"66",x"d4",x"87"),
  1432 => (x"a6",x"d8",x"80",x"c1"),
  1433 => (x"87",x"e7",x"c5",x"58"),
  1434 => (x"c1",x"48",x"66",x"d8"),
  1435 => (x"58",x"a6",x"dc",x"88"),
  1436 => (x"ff",x"87",x"dc",x"c5"),
  1437 => (x"70",x"87",x"f5",x"d8"),
  1438 => (x"87",x"d3",x"c5",x"4d"),
  1439 => (x"c0",x"48",x"66",x"cc"),
  1440 => (x"05",x"a8",x"66",x"e4"),
  1441 => (x"c0",x"87",x"f4",x"c4"),
  1442 => (x"c0",x"48",x"a6",x"e8"),
  1443 => (x"da",x"da",x"ff",x"78"),
  1444 => (x"ff",x"7e",x"70",x"87"),
  1445 => (x"c0",x"87",x"d4",x"da"),
  1446 => (x"c0",x"58",x"a6",x"f0"),
  1447 => (x"c0",x"05",x"a8",x"ec"),
  1448 => (x"48",x"a6",x"87",x"c7"),
  1449 => (x"c4",x"c0",x"78",x"6e"),
  1450 => (x"d7",x"d7",x"ff",x"87"),
  1451 => (x"49",x"66",x"d4",x"87"),
  1452 => (x"c4",x"c1",x"91",x"cc"),
  1453 => (x"80",x"71",x"48",x"66"),
  1454 => (x"c4",x"58",x"a6",x"c8"),
  1455 => (x"82",x"c8",x"4a",x"66"),
  1456 => (x"ca",x"49",x"66",x"c4"),
  1457 => (x"c0",x"51",x"6e",x"81"),
  1458 => (x"c1",x"49",x"66",x"ec"),
  1459 => (x"c1",x"89",x"6e",x"81"),
  1460 => (x"70",x"30",x"71",x"48"),
  1461 => (x"71",x"89",x"c1",x"49"),
  1462 => (x"e1",x"c2",x"7a",x"97"),
  1463 => (x"6e",x"49",x"bf",x"ec"),
  1464 => (x"4a",x"6a",x"97",x"29"),
  1465 => (x"c0",x"98",x"71",x"48"),
  1466 => (x"c4",x"58",x"a6",x"f4"),
  1467 => (x"80",x"c4",x"48",x"66"),
  1468 => (x"c8",x"58",x"a6",x"cc"),
  1469 => (x"c0",x"4c",x"bf",x"66"),
  1470 => (x"cc",x"48",x"66",x"e4"),
  1471 => (x"c0",x"02",x"a8",x"66"),
  1472 => (x"7e",x"c0",x"87",x"c5"),
  1473 => (x"c1",x"87",x"c2",x"c0"),
  1474 => (x"c0",x"1e",x"6e",x"7e"),
  1475 => (x"49",x"74",x"1e",x"e0"),
  1476 => (x"87",x"ec",x"d6",x"ff"),
  1477 => (x"4d",x"70",x"86",x"c8"),
  1478 => (x"06",x"ad",x"b7",x"c0"),
  1479 => (x"75",x"87",x"d4",x"c1"),
  1480 => (x"bf",x"66",x"c8",x"84"),
  1481 => (x"81",x"e0",x"c0",x"49"),
  1482 => (x"c1",x"4b",x"89",x"74"),
  1483 => (x"71",x"4a",x"dc",x"c1"),
  1484 => (x"87",x"ef",x"e7",x"fe"),
  1485 => (x"7e",x"74",x"84",x"c2"),
  1486 => (x"48",x"66",x"e8",x"c0"),
  1487 => (x"ec",x"c0",x"80",x"c1"),
  1488 => (x"f0",x"c0",x"58",x"a6"),
  1489 => (x"81",x"c1",x"49",x"66"),
  1490 => (x"c0",x"02",x"a9",x"70"),
  1491 => (x"4c",x"c0",x"87",x"c5"),
  1492 => (x"c1",x"87",x"c2",x"c0"),
  1493 => (x"cc",x"1e",x"74",x"4c"),
  1494 => (x"c0",x"49",x"bf",x"66"),
  1495 => (x"66",x"c4",x"81",x"e0"),
  1496 => (x"c8",x"1e",x"71",x"89"),
  1497 => (x"d5",x"ff",x"49",x"66"),
  1498 => (x"86",x"c8",x"87",x"d6"),
  1499 => (x"01",x"a8",x"b7",x"c0"),
  1500 => (x"c0",x"87",x"c5",x"ff"),
  1501 => (x"c0",x"02",x"66",x"e8"),
  1502 => (x"66",x"c4",x"87",x"d3"),
  1503 => (x"c0",x"81",x"c9",x"49"),
  1504 => (x"c4",x"51",x"66",x"e8"),
  1505 => (x"cd",x"c1",x"48",x"66"),
  1506 => (x"ce",x"c0",x"78",x"de"),
  1507 => (x"49",x"66",x"c4",x"87"),
  1508 => (x"51",x"c2",x"81",x"c9"),
  1509 => (x"c1",x"48",x"66",x"c4"),
  1510 => (x"d4",x"78",x"dc",x"cf"),
  1511 => (x"66",x"d8",x"48",x"66"),
  1512 => (x"cb",x"c0",x"04",x"a8"),
  1513 => (x"48",x"66",x"d4",x"87"),
  1514 => (x"a6",x"d8",x"80",x"c1"),
  1515 => (x"87",x"d1",x"c0",x"58"),
  1516 => (x"c1",x"48",x"66",x"d8"),
  1517 => (x"58",x"a6",x"dc",x"88"),
  1518 => (x"ff",x"87",x"c6",x"c0"),
  1519 => (x"70",x"87",x"ed",x"d3"),
  1520 => (x"48",x"a6",x"cc",x"4d"),
  1521 => (x"c6",x"c0",x"78",x"c0"),
  1522 => (x"df",x"d3",x"ff",x"87"),
  1523 => (x"c0",x"4d",x"70",x"87"),
  1524 => (x"c1",x"48",x"66",x"e0"),
  1525 => (x"a6",x"e4",x"c0",x"80"),
  1526 => (x"02",x"9d",x"75",x"58"),
  1527 => (x"d4",x"87",x"cb",x"c0"),
  1528 => (x"cc",x"c1",x"48",x"66"),
  1529 => (x"f4",x"04",x"a8",x"66"),
  1530 => (x"66",x"d4",x"87",x"da"),
  1531 => (x"03",x"a8",x"c7",x"48"),
  1532 => (x"d4",x"87",x"e1",x"c0"),
  1533 => (x"e2",x"c2",x"4c",x"66"),
  1534 => (x"78",x"c0",x"48",x"d0"),
  1535 => (x"91",x"cc",x"49",x"74"),
  1536 => (x"81",x"66",x"c4",x"c1"),
  1537 => (x"6a",x"4a",x"a1",x"c4"),
  1538 => (x"79",x"52",x"c0",x"4a"),
  1539 => (x"ac",x"c7",x"84",x"c1"),
  1540 => (x"87",x"e2",x"ff",x"04"),
  1541 => (x"02",x"66",x"e4",x"c0"),
  1542 => (x"c1",x"87",x"e2",x"c0"),
  1543 => (x"c1",x"49",x"66",x"c4"),
  1544 => (x"c4",x"c1",x"81",x"d4"),
  1545 => (x"dc",x"c1",x"4a",x"66"),
  1546 => (x"c1",x"52",x"c0",x"82"),
  1547 => (x"c1",x"79",x"d0",x"cc"),
  1548 => (x"c1",x"49",x"66",x"c4"),
  1549 => (x"c1",x"c1",x"81",x"d8"),
  1550 => (x"d6",x"c0",x"79",x"e0"),
  1551 => (x"66",x"c4",x"c1",x"87"),
  1552 => (x"81",x"d4",x"c1",x"49"),
  1553 => (x"4a",x"66",x"c4",x"c1"),
  1554 => (x"c1",x"82",x"d8",x"c1"),
  1555 => (x"c1",x"7a",x"e8",x"c1"),
  1556 => (x"c1",x"79",x"c7",x"cc"),
  1557 => (x"c1",x"49",x"66",x"c4"),
  1558 => (x"cf",x"c1",x"81",x"e0"),
  1559 => (x"d1",x"ff",x"79",x"ee"),
  1560 => (x"66",x"d0",x"87",x"c1"),
  1561 => (x"8e",x"cc",x"ff",x"48"),
  1562 => (x"4c",x"26",x"4d",x"26"),
  1563 => (x"4f",x"26",x"4b",x"26"),
  1564 => (x"c2",x"1e",x"c7",x"1e"),
  1565 => (x"1e",x"bf",x"cc",x"e2"),
  1566 => (x"1e",x"e4",x"e4",x"c1"),
  1567 => (x"97",x"f0",x"e1",x"c2"),
  1568 => (x"fb",x"ee",x"49",x"bf"),
  1569 => (x"e4",x"e4",x"c1",x"87"),
  1570 => (x"d9",x"e1",x"c0",x"49"),
  1571 => (x"26",x"8e",x"f4",x"87"),
  1572 => (x"e4",x"c1",x"1e",x"4f"),
  1573 => (x"50",x"c0",x"48",x"d8"),
  1574 => (x"bf",x"e0",x"d3",x"c2"),
  1575 => (x"f9",x"d5",x"ff",x"49"),
  1576 => (x"26",x"48",x"c0",x"87"),
  1577 => (x"1e",x"73",x"1e",x"4f"),
  1578 => (x"c2",x"87",x"c7",x"c7"),
  1579 => (x"c0",x"48",x"d8",x"e2"),
  1580 => (x"48",x"d4",x"ff",x"50"),
  1581 => (x"c1",x"78",x"ff",x"c3"),
  1582 => (x"fe",x"49",x"f0",x"c1"),
  1583 => (x"fe",x"87",x"e8",x"df"),
  1584 => (x"70",x"87",x"fd",x"ea"),
  1585 => (x"87",x"cd",x"02",x"98"),
  1586 => (x"87",x"f0",x"f2",x"fe"),
  1587 => (x"c4",x"02",x"98",x"70"),
  1588 => (x"c2",x"4a",x"c1",x"87"),
  1589 => (x"72",x"4a",x"c0",x"87"),
  1590 => (x"87",x"c8",x"02",x"9a"),
  1591 => (x"49",x"fc",x"c1",x"c1"),
  1592 => (x"87",x"c3",x"df",x"fe"),
  1593 => (x"48",x"cc",x"e2",x"c2"),
  1594 => (x"e1",x"c2",x"78",x"c0"),
  1595 => (x"50",x"c0",x"48",x"f0"),
  1596 => (x"87",x"fc",x"fd",x"49"),
  1597 => (x"70",x"87",x"da",x"fe"),
  1598 => (x"ce",x"02",x"9b",x"4b"),
  1599 => (x"c0",x"e6",x"c1",x"87"),
  1600 => (x"de",x"49",x"c7",x"5b"),
  1601 => (x"49",x"c1",x"87",x"d2"),
  1602 => (x"c2",x"87",x"ee",x"df"),
  1603 => (x"e1",x"c0",x"87",x"ed"),
  1604 => (x"87",x"fa",x"87",x"cf"),
  1605 => (x"4f",x"26",x"4b",x"26"),
  1606 => (x"00",x"00",x"00",x"00"),
  1607 => (x"00",x"00",x"00",x"00"),
  1608 => (x"00",x"00",x"00",x"01"),
  1609 => (x"00",x"00",x"0f",x"ba"),
  1610 => (x"00",x"00",x"28",x"a4"),
  1611 => (x"00",x"00",x"00",x"00"),
  1612 => (x"00",x"00",x"0f",x"ba"),
  1613 => (x"00",x"00",x"28",x"c2"),
  1614 => (x"00",x"00",x"00",x"00"),
  1615 => (x"00",x"00",x"0f",x"ba"),
  1616 => (x"00",x"00",x"28",x"e0"),
  1617 => (x"00",x"00",x"00",x"00"),
  1618 => (x"00",x"00",x"0f",x"ba"),
  1619 => (x"00",x"00",x"28",x"fe"),
  1620 => (x"00",x"00",x"00",x"00"),
  1621 => (x"00",x"00",x"0f",x"ba"),
  1622 => (x"00",x"00",x"29",x"1c"),
  1623 => (x"00",x"00",x"00",x"00"),
  1624 => (x"00",x"00",x"0f",x"ba"),
  1625 => (x"00",x"00",x"29",x"3a"),
  1626 => (x"00",x"00",x"00",x"00"),
  1627 => (x"00",x"00",x"0f",x"ba"),
  1628 => (x"00",x"00",x"29",x"58"),
  1629 => (x"00",x"00",x"00",x"00"),
  1630 => (x"00",x"00",x"13",x"10"),
  1631 => (x"00",x"00",x"00",x"00"),
  1632 => (x"00",x"00",x"00",x"00"),
  1633 => (x"00",x"00",x"10",x"b4"),
  1634 => (x"00",x"00",x"00",x"00"),
  1635 => (x"00",x"00",x"00",x"00"),
  1636 => (x"00",x"00",x"10",x"80"),
  1637 => (x"db",x"86",x"fc",x"1e"),
  1638 => (x"fc",x"7e",x"70",x"87"),
  1639 => (x"1e",x"4f",x"26",x"8e"),
  1640 => (x"c0",x"48",x"f0",x"fe"),
  1641 => (x"79",x"09",x"cd",x"78"),
  1642 => (x"1e",x"4f",x"26",x"09"),
  1643 => (x"49",x"d4",x"e6",x"c1"),
  1644 => (x"4f",x"26",x"87",x"ed"),
  1645 => (x"bf",x"f0",x"fe",x"1e"),
  1646 => (x"1e",x"4f",x"26",x"48"),
  1647 => (x"c1",x"48",x"f0",x"fe"),
  1648 => (x"1e",x"4f",x"26",x"78"),
  1649 => (x"c0",x"48",x"f0",x"fe"),
  1650 => (x"1e",x"4f",x"26",x"78"),
  1651 => (x"52",x"c0",x"4a",x"71"),
  1652 => (x"0e",x"4f",x"26",x"51"),
  1653 => (x"5d",x"5c",x"5b",x"5e"),
  1654 => (x"71",x"86",x"f4",x"0e"),
  1655 => (x"7e",x"6d",x"97",x"4d"),
  1656 => (x"97",x"4c",x"a5",x"c1"),
  1657 => (x"a6",x"c8",x"48",x"6c"),
  1658 => (x"c4",x"48",x"6e",x"58"),
  1659 => (x"c5",x"05",x"a8",x"66"),
  1660 => (x"c0",x"48",x"ff",x"87"),
  1661 => (x"ca",x"ff",x"87",x"e6"),
  1662 => (x"49",x"a5",x"c2",x"87"),
  1663 => (x"71",x"4b",x"6c",x"97"),
  1664 => (x"6b",x"97",x"4b",x"a3"),
  1665 => (x"7e",x"6c",x"97",x"4b"),
  1666 => (x"80",x"c1",x"48",x"6e"),
  1667 => (x"c7",x"58",x"a6",x"c8"),
  1668 => (x"58",x"a6",x"cc",x"98"),
  1669 => (x"fe",x"7c",x"97",x"70"),
  1670 => (x"48",x"73",x"87",x"e1"),
  1671 => (x"4d",x"26",x"8e",x"f4"),
  1672 => (x"4b",x"26",x"4c",x"26"),
  1673 => (x"73",x"1e",x"4f",x"26"),
  1674 => (x"fe",x"86",x"f4",x"1e"),
  1675 => (x"bf",x"e0",x"87",x"d5"),
  1676 => (x"e0",x"c0",x"49",x"4b"),
  1677 => (x"c0",x"02",x"99",x"c0"),
  1678 => (x"4a",x"73",x"87",x"ea"),
  1679 => (x"c2",x"9a",x"ff",x"c3"),
  1680 => (x"bf",x"97",x"cc",x"e6"),
  1681 => (x"ce",x"e6",x"c2",x"49"),
  1682 => (x"c2",x"51",x"72",x"81"),
  1683 => (x"bf",x"97",x"cc",x"e6"),
  1684 => (x"c1",x"48",x"6e",x"7e"),
  1685 => (x"58",x"a6",x"c8",x"80"),
  1686 => (x"a6",x"cc",x"98",x"c7"),
  1687 => (x"cc",x"e6",x"c2",x"58"),
  1688 => (x"50",x"66",x"c8",x"48"),
  1689 => (x"70",x"87",x"cd",x"fd"),
  1690 => (x"87",x"cf",x"fd",x"7e"),
  1691 => (x"4b",x"26",x"8e",x"f4"),
  1692 => (x"c2",x"1e",x"4f",x"26"),
  1693 => (x"fd",x"49",x"cc",x"e6"),
  1694 => (x"e8",x"c1",x"87",x"d1"),
  1695 => (x"de",x"fc",x"49",x"e6"),
  1696 => (x"87",x"e8",x"c4",x"87"),
  1697 => (x"5e",x"0e",x"4f",x"26"),
  1698 => (x"0e",x"5d",x"5c",x"5b"),
  1699 => (x"7e",x"71",x"86",x"fc"),
  1700 => (x"c2",x"4d",x"d4",x"ff"),
  1701 => (x"fc",x"49",x"cc",x"e6"),
  1702 => (x"4b",x"70",x"87",x"f9"),
  1703 => (x"04",x"ab",x"b7",x"c0"),
  1704 => (x"c3",x"87",x"f5",x"c2"),
  1705 => (x"c9",x"05",x"ab",x"f0"),
  1706 => (x"e4",x"ed",x"c1",x"87"),
  1707 => (x"c2",x"78",x"c1",x"48"),
  1708 => (x"e0",x"c3",x"87",x"d6"),
  1709 => (x"87",x"c9",x"05",x"ab"),
  1710 => (x"48",x"e8",x"ed",x"c1"),
  1711 => (x"c7",x"c2",x"78",x"c1"),
  1712 => (x"e8",x"ed",x"c1",x"87"),
  1713 => (x"87",x"c6",x"02",x"bf"),
  1714 => (x"4c",x"a3",x"c0",x"c2"),
  1715 => (x"4c",x"73",x"87",x"c2"),
  1716 => (x"bf",x"e4",x"ed",x"c1"),
  1717 => (x"87",x"e0",x"c0",x"02"),
  1718 => (x"b7",x"c4",x"49",x"74"),
  1719 => (x"ed",x"c1",x"91",x"29"),
  1720 => (x"4a",x"74",x"81",x"ec"),
  1721 => (x"92",x"c2",x"9a",x"cf"),
  1722 => (x"30",x"72",x"48",x"c1"),
  1723 => (x"ba",x"ff",x"4a",x"70"),
  1724 => (x"98",x"69",x"48",x"72"),
  1725 => (x"87",x"db",x"79",x"70"),
  1726 => (x"b7",x"c4",x"49",x"74"),
  1727 => (x"ed",x"c1",x"91",x"29"),
  1728 => (x"4a",x"74",x"81",x"ec"),
  1729 => (x"92",x"c2",x"9a",x"cf"),
  1730 => (x"30",x"72",x"48",x"c3"),
  1731 => (x"69",x"48",x"4a",x"70"),
  1732 => (x"6e",x"79",x"70",x"b0"),
  1733 => (x"87",x"e4",x"c0",x"05"),
  1734 => (x"c8",x"48",x"d0",x"ff"),
  1735 => (x"7d",x"c5",x"78",x"e1"),
  1736 => (x"bf",x"e8",x"ed",x"c1"),
  1737 => (x"c3",x"87",x"c3",x"02"),
  1738 => (x"ed",x"c1",x"7d",x"e0"),
  1739 => (x"c3",x"02",x"bf",x"e4"),
  1740 => (x"7d",x"f0",x"c3",x"87"),
  1741 => (x"d0",x"ff",x"7d",x"73"),
  1742 => (x"78",x"e0",x"c0",x"48"),
  1743 => (x"48",x"e8",x"ed",x"c1"),
  1744 => (x"ed",x"c1",x"78",x"c0"),
  1745 => (x"78",x"c0",x"48",x"e4"),
  1746 => (x"49",x"cc",x"e6",x"c2"),
  1747 => (x"70",x"87",x"c4",x"fa"),
  1748 => (x"ab",x"b7",x"c0",x"4b"),
  1749 => (x"87",x"cb",x"fd",x"03"),
  1750 => (x"8e",x"fc",x"48",x"c0"),
  1751 => (x"4c",x"26",x"4d",x"26"),
  1752 => (x"4f",x"26",x"4b",x"26"),
  1753 => (x"00",x"00",x"00",x"00"),
  1754 => (x"00",x"00",x"00",x"00"),
  1755 => (x"00",x"00",x"00",x"00"),
  1756 => (x"00",x"00",x"00",x"00"),
  1757 => (x"00",x"00",x"00",x"00"),
  1758 => (x"00",x"00",x"00",x"00"),
  1759 => (x"00",x"00",x"00",x"00"),
  1760 => (x"00",x"00",x"00",x"00"),
  1761 => (x"00",x"00",x"00",x"00"),
  1762 => (x"00",x"00",x"00",x"00"),
  1763 => (x"00",x"00",x"00",x"00"),
  1764 => (x"00",x"00",x"00",x"00"),
  1765 => (x"00",x"00",x"00",x"00"),
  1766 => (x"00",x"00",x"00",x"00"),
  1767 => (x"00",x"00",x"00",x"00"),
  1768 => (x"00",x"00",x"00",x"00"),
  1769 => (x"00",x"00",x"00",x"00"),
  1770 => (x"00",x"00",x"00",x"00"),
  1771 => (x"72",x"4a",x"c0",x"1e"),
  1772 => (x"c1",x"91",x"c4",x"49"),
  1773 => (x"c0",x"81",x"ec",x"ed"),
  1774 => (x"d0",x"82",x"c1",x"79"),
  1775 => (x"ee",x"04",x"aa",x"b7"),
  1776 => (x"0e",x"4f",x"26",x"87"),
  1777 => (x"5d",x"5c",x"5b",x"5e"),
  1778 => (x"f7",x"4d",x"71",x"0e"),
  1779 => (x"4a",x"75",x"87",x"f5"),
  1780 => (x"92",x"2a",x"b7",x"c4"),
  1781 => (x"82",x"ec",x"ed",x"c1"),
  1782 => (x"9c",x"cf",x"4c",x"75"),
  1783 => (x"49",x"6a",x"94",x"c2"),
  1784 => (x"c3",x"2b",x"74",x"4b"),
  1785 => (x"74",x"48",x"c2",x"9b"),
  1786 => (x"ff",x"4c",x"70",x"30"),
  1787 => (x"71",x"48",x"74",x"bc"),
  1788 => (x"f7",x"7a",x"70",x"98"),
  1789 => (x"48",x"73",x"87",x"c5"),
  1790 => (x"4c",x"26",x"4d",x"26"),
  1791 => (x"4f",x"26",x"4b",x"26"),
  1792 => (x"48",x"d0",x"ff",x"1e"),
  1793 => (x"71",x"78",x"e1",x"c8"),
  1794 => (x"08",x"d4",x"ff",x"48"),
  1795 => (x"48",x"66",x"c4",x"78"),
  1796 => (x"78",x"08",x"d4",x"ff"),
  1797 => (x"71",x"1e",x"4f",x"26"),
  1798 => (x"49",x"66",x"c4",x"4a"),
  1799 => (x"ff",x"49",x"72",x"1e"),
  1800 => (x"d0",x"ff",x"87",x"de"),
  1801 => (x"78",x"e0",x"c0",x"48"),
  1802 => (x"4f",x"26",x"8e",x"fc"),
  1803 => (x"71",x"1e",x"73",x"1e"),
  1804 => (x"49",x"66",x"c8",x"4b"),
  1805 => (x"c1",x"4a",x"73",x"1e"),
  1806 => (x"ff",x"49",x"a2",x"e0"),
  1807 => (x"8e",x"fc",x"87",x"d8"),
  1808 => (x"4f",x"26",x"4b",x"26"),
  1809 => (x"48",x"d0",x"ff",x"1e"),
  1810 => (x"71",x"78",x"c9",x"c8"),
  1811 => (x"08",x"d4",x"ff",x"48"),
  1812 => (x"1e",x"4f",x"26",x"78"),
  1813 => (x"eb",x"49",x"4a",x"71"),
  1814 => (x"48",x"d0",x"ff",x"87"),
  1815 => (x"4f",x"26",x"78",x"c8"),
  1816 => (x"71",x"1e",x"73",x"1e"),
  1817 => (x"e4",x"e6",x"c2",x"4b"),
  1818 => (x"87",x"c3",x"02",x"bf"),
  1819 => (x"ff",x"87",x"eb",x"c2"),
  1820 => (x"c9",x"c8",x"48",x"d0"),
  1821 => (x"c0",x"48",x"73",x"78"),
  1822 => (x"d4",x"ff",x"b0",x"e0"),
  1823 => (x"e6",x"c2",x"78",x"08"),
  1824 => (x"78",x"c0",x"48",x"d8"),
  1825 => (x"c5",x"02",x"66",x"c8"),
  1826 => (x"49",x"ff",x"c3",x"87"),
  1827 => (x"49",x"c0",x"87",x"c2"),
  1828 => (x"59",x"e0",x"e6",x"c2"),
  1829 => (x"c6",x"02",x"66",x"cc"),
  1830 => (x"d5",x"d5",x"c5",x"87"),
  1831 => (x"cf",x"87",x"c4",x"4a"),
  1832 => (x"c2",x"4a",x"ff",x"ff"),
  1833 => (x"c2",x"5a",x"e4",x"e6"),
  1834 => (x"c1",x"48",x"e4",x"e6"),
  1835 => (x"26",x"4b",x"26",x"78"),
  1836 => (x"5b",x"5e",x"0e",x"4f"),
  1837 => (x"71",x"0e",x"5d",x"5c"),
  1838 => (x"e0",x"e6",x"c2",x"4d"),
  1839 => (x"9d",x"75",x"4b",x"bf"),
  1840 => (x"49",x"87",x"cb",x"02"),
  1841 => (x"f1",x"c1",x"91",x"c8"),
  1842 => (x"82",x"71",x"4a",x"d8"),
  1843 => (x"f5",x"c1",x"87",x"c4"),
  1844 => (x"4c",x"c0",x"4a",x"d8"),
  1845 => (x"99",x"73",x"49",x"12"),
  1846 => (x"bf",x"dc",x"e6",x"c2"),
  1847 => (x"ff",x"b8",x"71",x"48"),
  1848 => (x"c1",x"78",x"08",x"d4"),
  1849 => (x"c8",x"84",x"2b",x"b7"),
  1850 => (x"e7",x"04",x"ac",x"b7"),
  1851 => (x"d8",x"e6",x"c2",x"87"),
  1852 => (x"80",x"c8",x"48",x"bf"),
  1853 => (x"58",x"dc",x"e6",x"c2"),
  1854 => (x"4c",x"26",x"4d",x"26"),
  1855 => (x"4f",x"26",x"4b",x"26"),
  1856 => (x"71",x"1e",x"73",x"1e"),
  1857 => (x"9a",x"4a",x"13",x"4b"),
  1858 => (x"72",x"87",x"cb",x"02"),
  1859 => (x"87",x"e1",x"fe",x"49"),
  1860 => (x"05",x"9a",x"4a",x"13"),
  1861 => (x"4b",x"26",x"87",x"f5"),
  1862 => (x"c2",x"1e",x"4f",x"26"),
  1863 => (x"49",x"bf",x"d8",x"e6"),
  1864 => (x"48",x"d8",x"e6",x"c2"),
  1865 => (x"c4",x"78",x"a1",x"c1"),
  1866 => (x"03",x"a9",x"b7",x"c0"),
  1867 => (x"d4",x"ff",x"87",x"db"),
  1868 => (x"dc",x"e6",x"c2",x"48"),
  1869 => (x"e6",x"c2",x"78",x"bf"),
  1870 => (x"c2",x"49",x"bf",x"d8"),
  1871 => (x"c1",x"48",x"d8",x"e6"),
  1872 => (x"c0",x"c4",x"78",x"a1"),
  1873 => (x"e5",x"04",x"a9",x"b7"),
  1874 => (x"48",x"d0",x"ff",x"87"),
  1875 => (x"e6",x"c2",x"78",x"c8"),
  1876 => (x"78",x"c0",x"48",x"e4"),
  1877 => (x"00",x"00",x"4f",x"26"),
  1878 => (x"00",x"00",x"00",x"00"),
  1879 => (x"00",x"00",x"00",x"00"),
  1880 => (x"5f",x"00",x"00",x"00"),
  1881 => (x"00",x"00",x"00",x"5f"),
  1882 => (x"00",x"03",x"03",x"00"),
  1883 => (x"00",x"00",x"03",x"03"),
  1884 => (x"14",x"7f",x"7f",x"14"),
  1885 => (x"00",x"14",x"7f",x"7f"),
  1886 => (x"6b",x"2e",x"24",x"00"),
  1887 => (x"00",x"12",x"3a",x"6b"),
  1888 => (x"18",x"36",x"6a",x"4c"),
  1889 => (x"00",x"32",x"56",x"6c"),
  1890 => (x"59",x"4f",x"7e",x"30"),
  1891 => (x"40",x"68",x"3a",x"77"),
  1892 => (x"07",x"04",x"00",x"00"),
  1893 => (x"00",x"00",x"00",x"03"),
  1894 => (x"3e",x"1c",x"00",x"00"),
  1895 => (x"00",x"00",x"41",x"63"),
  1896 => (x"63",x"41",x"00",x"00"),
  1897 => (x"00",x"00",x"1c",x"3e"),
  1898 => (x"1c",x"3e",x"2a",x"08"),
  1899 => (x"08",x"2a",x"3e",x"1c"),
  1900 => (x"3e",x"08",x"08",x"00"),
  1901 => (x"00",x"08",x"08",x"3e"),
  1902 => (x"e0",x"80",x"00",x"00"),
  1903 => (x"00",x"00",x"00",x"60"),
  1904 => (x"08",x"08",x"08",x"00"),
  1905 => (x"00",x"08",x"08",x"08"),
  1906 => (x"60",x"00",x"00",x"00"),
  1907 => (x"00",x"00",x"00",x"60"),
  1908 => (x"18",x"30",x"60",x"40"),
  1909 => (x"01",x"03",x"06",x"0c"),
  1910 => (x"59",x"7f",x"3e",x"00"),
  1911 => (x"00",x"3e",x"7f",x"4d"),
  1912 => (x"7f",x"06",x"04",x"00"),
  1913 => (x"00",x"00",x"00",x"7f"),
  1914 => (x"71",x"63",x"42",x"00"),
  1915 => (x"00",x"46",x"4f",x"59"),
  1916 => (x"49",x"63",x"22",x"00"),
  1917 => (x"00",x"36",x"7f",x"49"),
  1918 => (x"13",x"16",x"1c",x"18"),
  1919 => (x"00",x"10",x"7f",x"7f"),
  1920 => (x"45",x"67",x"27",x"00"),
  1921 => (x"00",x"39",x"7d",x"45"),
  1922 => (x"4b",x"7e",x"3c",x"00"),
  1923 => (x"00",x"30",x"79",x"49"),
  1924 => (x"71",x"01",x"01",x"00"),
  1925 => (x"00",x"07",x"0f",x"79"),
  1926 => (x"49",x"7f",x"36",x"00"),
  1927 => (x"00",x"36",x"7f",x"49"),
  1928 => (x"49",x"4f",x"06",x"00"),
  1929 => (x"00",x"1e",x"3f",x"69"),
  1930 => (x"66",x"00",x"00",x"00"),
  1931 => (x"00",x"00",x"00",x"66"),
  1932 => (x"e6",x"80",x"00",x"00"),
  1933 => (x"00",x"00",x"00",x"66"),
  1934 => (x"14",x"08",x"08",x"00"),
  1935 => (x"00",x"22",x"22",x"14"),
  1936 => (x"14",x"14",x"14",x"00"),
  1937 => (x"00",x"14",x"14",x"14"),
  1938 => (x"14",x"22",x"22",x"00"),
  1939 => (x"00",x"08",x"08",x"14"),
  1940 => (x"51",x"03",x"02",x"00"),
  1941 => (x"00",x"06",x"0f",x"59"),
  1942 => (x"5d",x"41",x"7f",x"3e"),
  1943 => (x"00",x"1e",x"1f",x"55"),
  1944 => (x"09",x"7f",x"7e",x"00"),
  1945 => (x"00",x"7e",x"7f",x"09"),
  1946 => (x"49",x"7f",x"7f",x"00"),
  1947 => (x"00",x"36",x"7f",x"49"),
  1948 => (x"63",x"3e",x"1c",x"00"),
  1949 => (x"00",x"41",x"41",x"41"),
  1950 => (x"41",x"7f",x"7f",x"00"),
  1951 => (x"00",x"1c",x"3e",x"63"),
  1952 => (x"49",x"7f",x"7f",x"00"),
  1953 => (x"00",x"41",x"41",x"49"),
  1954 => (x"09",x"7f",x"7f",x"00"),
  1955 => (x"00",x"01",x"01",x"09"),
  1956 => (x"41",x"7f",x"3e",x"00"),
  1957 => (x"00",x"7a",x"7b",x"49"),
  1958 => (x"08",x"7f",x"7f",x"00"),
  1959 => (x"00",x"7f",x"7f",x"08"),
  1960 => (x"7f",x"41",x"00",x"00"),
  1961 => (x"00",x"00",x"41",x"7f"),
  1962 => (x"40",x"60",x"20",x"00"),
  1963 => (x"00",x"3f",x"7f",x"40"),
  1964 => (x"1c",x"08",x"7f",x"7f"),
  1965 => (x"00",x"41",x"63",x"36"),
  1966 => (x"40",x"7f",x"7f",x"00"),
  1967 => (x"00",x"40",x"40",x"40"),
  1968 => (x"0c",x"06",x"7f",x"7f"),
  1969 => (x"00",x"7f",x"7f",x"06"),
  1970 => (x"0c",x"06",x"7f",x"7f"),
  1971 => (x"00",x"7f",x"7f",x"18"),
  1972 => (x"41",x"7f",x"3e",x"00"),
  1973 => (x"00",x"3e",x"7f",x"41"),
  1974 => (x"09",x"7f",x"7f",x"00"),
  1975 => (x"00",x"06",x"0f",x"09"),
  1976 => (x"61",x"41",x"7f",x"3e"),
  1977 => (x"00",x"40",x"7e",x"7f"),
  1978 => (x"09",x"7f",x"7f",x"00"),
  1979 => (x"00",x"66",x"7f",x"19"),
  1980 => (x"4d",x"6f",x"26",x"00"),
  1981 => (x"00",x"32",x"7b",x"59"),
  1982 => (x"7f",x"01",x"01",x"00"),
  1983 => (x"00",x"01",x"01",x"7f"),
  1984 => (x"40",x"7f",x"3f",x"00"),
  1985 => (x"00",x"3f",x"7f",x"40"),
  1986 => (x"70",x"3f",x"0f",x"00"),
  1987 => (x"00",x"0f",x"3f",x"70"),
  1988 => (x"18",x"30",x"7f",x"7f"),
  1989 => (x"00",x"7f",x"7f",x"30"),
  1990 => (x"1c",x"36",x"63",x"41"),
  1991 => (x"41",x"63",x"36",x"1c"),
  1992 => (x"7c",x"06",x"03",x"01"),
  1993 => (x"01",x"03",x"06",x"7c"),
  1994 => (x"4d",x"59",x"71",x"61"),
  1995 => (x"00",x"41",x"43",x"47"),
  1996 => (x"7f",x"7f",x"00",x"00"),
  1997 => (x"00",x"00",x"41",x"41"),
  1998 => (x"0c",x"06",x"03",x"01"),
  1999 => (x"40",x"60",x"30",x"18"),
  2000 => (x"41",x"41",x"00",x"00"),
  2001 => (x"00",x"00",x"7f",x"7f"),
  2002 => (x"03",x"06",x"0c",x"08"),
  2003 => (x"00",x"08",x"0c",x"06"),
  2004 => (x"80",x"80",x"80",x"80"),
  2005 => (x"00",x"80",x"80",x"80"),
  2006 => (x"03",x"00",x"00",x"00"),
  2007 => (x"00",x"00",x"04",x"07"),
  2008 => (x"54",x"74",x"20",x"00"),
  2009 => (x"00",x"78",x"7c",x"54"),
  2010 => (x"44",x"7f",x"7f",x"00"),
  2011 => (x"00",x"38",x"7c",x"44"),
  2012 => (x"44",x"7c",x"38",x"00"),
  2013 => (x"00",x"00",x"44",x"44"),
  2014 => (x"44",x"7c",x"38",x"00"),
  2015 => (x"00",x"7f",x"7f",x"44"),
  2016 => (x"54",x"7c",x"38",x"00"),
  2017 => (x"00",x"18",x"5c",x"54"),
  2018 => (x"7f",x"7e",x"04",x"00"),
  2019 => (x"00",x"00",x"05",x"05"),
  2020 => (x"a4",x"bc",x"18",x"00"),
  2021 => (x"00",x"7c",x"fc",x"a4"),
  2022 => (x"04",x"7f",x"7f",x"00"),
  2023 => (x"00",x"78",x"7c",x"04"),
  2024 => (x"3d",x"00",x"00",x"00"),
  2025 => (x"00",x"00",x"40",x"7d"),
  2026 => (x"80",x"80",x"80",x"00"),
  2027 => (x"00",x"00",x"7d",x"fd"),
  2028 => (x"10",x"7f",x"7f",x"00"),
  2029 => (x"00",x"44",x"6c",x"38"),
  2030 => (x"3f",x"00",x"00",x"00"),
  2031 => (x"00",x"00",x"40",x"7f"),
  2032 => (x"18",x"0c",x"7c",x"7c"),
  2033 => (x"00",x"78",x"7c",x"0c"),
  2034 => (x"04",x"7c",x"7c",x"00"),
  2035 => (x"00",x"78",x"7c",x"04"),
  2036 => (x"44",x"7c",x"38",x"00"),
  2037 => (x"00",x"38",x"7c",x"44"),
  2038 => (x"24",x"fc",x"fc",x"00"),
  2039 => (x"00",x"18",x"3c",x"24"),
  2040 => (x"24",x"3c",x"18",x"00"),
  2041 => (x"00",x"fc",x"fc",x"24"),
  2042 => (x"04",x"7c",x"7c",x"00"),
  2043 => (x"00",x"08",x"0c",x"04"),
  2044 => (x"54",x"5c",x"48",x"00"),
  2045 => (x"00",x"20",x"74",x"54"),
  2046 => (x"7f",x"3f",x"04",x"00"),
  2047 => (x"00",x"00",x"44",x"44"),
  2048 => (x"40",x"7c",x"3c",x"00"),
  2049 => (x"00",x"7c",x"7c",x"40"),
  2050 => (x"60",x"3c",x"1c",x"00"),
  2051 => (x"00",x"1c",x"3c",x"60"),
  2052 => (x"30",x"60",x"7c",x"3c"),
  2053 => (x"00",x"3c",x"7c",x"60"),
  2054 => (x"10",x"38",x"6c",x"44"),
  2055 => (x"00",x"44",x"6c",x"38"),
  2056 => (x"e0",x"bc",x"1c",x"00"),
  2057 => (x"00",x"1c",x"3c",x"60"),
  2058 => (x"74",x"64",x"44",x"00"),
  2059 => (x"00",x"44",x"4c",x"5c"),
  2060 => (x"3e",x"08",x"08",x"00"),
  2061 => (x"00",x"41",x"41",x"77"),
  2062 => (x"7f",x"00",x"00",x"00"),
  2063 => (x"00",x"00",x"00",x"7f"),
  2064 => (x"77",x"41",x"41",x"00"),
  2065 => (x"00",x"08",x"08",x"3e"),
  2066 => (x"03",x"01",x"01",x"02"),
  2067 => (x"00",x"01",x"02",x"02"),
  2068 => (x"7f",x"7f",x"7f",x"7f"),
  2069 => (x"00",x"7f",x"7f",x"7f"),
  2070 => (x"1c",x"1c",x"08",x"08"),
  2071 => (x"7f",x"7f",x"3e",x"3e"),
  2072 => (x"3e",x"3e",x"7f",x"7f"),
  2073 => (x"08",x"08",x"1c",x"1c"),
  2074 => (x"7c",x"18",x"10",x"00"),
  2075 => (x"00",x"10",x"18",x"7c"),
  2076 => (x"7c",x"30",x"10",x"00"),
  2077 => (x"00",x"10",x"30",x"7c"),
  2078 => (x"60",x"60",x"30",x"10"),
  2079 => (x"00",x"06",x"1e",x"78"),
  2080 => (x"18",x"3c",x"66",x"42"),
  2081 => (x"00",x"42",x"66",x"3c"),
  2082 => (x"c2",x"6a",x"38",x"78"),
  2083 => (x"00",x"38",x"6c",x"c6"),
  2084 => (x"60",x"00",x"00",x"60"),
  2085 => (x"00",x"60",x"00",x"00"),
  2086 => (x"5c",x"5b",x"5e",x"0e"),
  2087 => (x"86",x"fc",x"0e",x"5d"),
  2088 => (x"e6",x"c2",x"7e",x"71"),
  2089 => (x"c0",x"4c",x"bf",x"ec"),
  2090 => (x"c4",x"1e",x"c0",x"4b"),
  2091 => (x"c4",x"02",x"ab",x"66"),
  2092 => (x"c2",x"4d",x"c0",x"87"),
  2093 => (x"75",x"4d",x"c1",x"87"),
  2094 => (x"ee",x"49",x"73",x"1e"),
  2095 => (x"86",x"c8",x"87",x"e2"),
  2096 => (x"ef",x"49",x"e0",x"c0"),
  2097 => (x"a4",x"c4",x"87",x"eb"),
  2098 => (x"f0",x"49",x"6a",x"4a"),
  2099 => (x"c9",x"f1",x"87",x"f2"),
  2100 => (x"c1",x"84",x"cc",x"87"),
  2101 => (x"ab",x"b7",x"c8",x"83"),
  2102 => (x"87",x"cd",x"ff",x"04"),
  2103 => (x"4d",x"26",x"8e",x"fc"),
  2104 => (x"4b",x"26",x"4c",x"26"),
  2105 => (x"71",x"1e",x"4f",x"26"),
  2106 => (x"f0",x"e6",x"c2",x"4a"),
  2107 => (x"f0",x"e6",x"c2",x"5a"),
  2108 => (x"49",x"78",x"c7",x"48"),
  2109 => (x"26",x"87",x"e1",x"fe"),
  2110 => (x"1e",x"73",x"1e",x"4f"),
  2111 => (x"b7",x"c0",x"4a",x"71"),
  2112 => (x"87",x"d3",x"03",x"aa"),
  2113 => (x"bf",x"e4",x"d2",x"c2"),
  2114 => (x"c1",x"87",x"c4",x"05"),
  2115 => (x"c0",x"87",x"c2",x"4b"),
  2116 => (x"e8",x"d2",x"c2",x"4b"),
  2117 => (x"c2",x"87",x"c4",x"5b"),
  2118 => (x"fc",x"5a",x"e8",x"d2"),
  2119 => (x"e4",x"d2",x"c2",x"48"),
  2120 => (x"c1",x"4a",x"78",x"bf"),
  2121 => (x"a2",x"c0",x"c1",x"9a"),
  2122 => (x"87",x"e7",x"ec",x"49"),
  2123 => (x"4f",x"26",x"4b",x"26"),
  2124 => (x"c4",x"4a",x"71",x"1e"),
  2125 => (x"49",x"72",x"1e",x"66"),
  2126 => (x"fc",x"87",x"f1",x"eb"),
  2127 => (x"1e",x"4f",x"26",x"8e"),
  2128 => (x"c3",x"48",x"d4",x"ff"),
  2129 => (x"d0",x"ff",x"78",x"ff"),
  2130 => (x"78",x"e1",x"c0",x"48"),
  2131 => (x"c1",x"48",x"d4",x"ff"),
  2132 => (x"c4",x"48",x"71",x"78"),
  2133 => (x"08",x"d4",x"ff",x"30"),
  2134 => (x"48",x"d0",x"ff",x"78"),
  2135 => (x"26",x"78",x"e0",x"c0"),
  2136 => (x"5b",x"5e",x"0e",x"4f"),
  2137 => (x"f0",x"0e",x"5d",x"5c"),
  2138 => (x"c8",x"7e",x"c0",x"86"),
  2139 => (x"bf",x"ec",x"48",x"a6"),
  2140 => (x"c2",x"80",x"fc",x"78"),
  2141 => (x"78",x"bf",x"ec",x"e6"),
  2142 => (x"bf",x"f4",x"e6",x"c2"),
  2143 => (x"4c",x"bf",x"e8",x"4d"),
  2144 => (x"bf",x"e4",x"d2",x"c2"),
  2145 => (x"87",x"fe",x"e3",x"49"),
  2146 => (x"f6",x"e8",x"49",x"c7"),
  2147 => (x"c2",x"49",x"70",x"87"),
  2148 => (x"87",x"d0",x"05",x"99"),
  2149 => (x"bf",x"dc",x"d2",x"c2"),
  2150 => (x"c8",x"b9",x"ff",x"49"),
  2151 => (x"99",x"c1",x"99",x"66"),
  2152 => (x"87",x"c2",x"c2",x"02"),
  2153 => (x"cb",x"49",x"e8",x"cf"),
  2154 => (x"a6",x"d0",x"87",x"fe"),
  2155 => (x"e8",x"49",x"c7",x"58"),
  2156 => (x"98",x"70",x"87",x"d1"),
  2157 => (x"c8",x"87",x"c9",x"05"),
  2158 => (x"99",x"c1",x"49",x"66"),
  2159 => (x"87",x"c6",x"c1",x"02"),
  2160 => (x"c8",x"4b",x"66",x"cc"),
  2161 => (x"bf",x"ec",x"48",x"a6"),
  2162 => (x"e4",x"d2",x"c2",x"78"),
  2163 => (x"f5",x"e2",x"49",x"bf"),
  2164 => (x"cb",x"49",x"73",x"87"),
  2165 => (x"98",x"70",x"87",x"de"),
  2166 => (x"c2",x"87",x"d7",x"02"),
  2167 => (x"49",x"bf",x"d8",x"d2"),
  2168 => (x"d2",x"c2",x"b9",x"c1"),
  2169 => (x"fd",x"71",x"59",x"dc"),
  2170 => (x"e8",x"cf",x"87",x"d5"),
  2171 => (x"87",x"f8",x"ca",x"49"),
  2172 => (x"49",x"c7",x"4b",x"70"),
  2173 => (x"70",x"87",x"cc",x"e7"),
  2174 => (x"c6",x"ff",x"05",x"98"),
  2175 => (x"49",x"66",x"c8",x"87"),
  2176 => (x"fe",x"05",x"99",x"c1"),
  2177 => (x"d2",x"c2",x"87",x"fd"),
  2178 => (x"c1",x"4a",x"bf",x"e4"),
  2179 => (x"e8",x"d2",x"c2",x"ba"),
  2180 => (x"7a",x"0a",x"fc",x"5a"),
  2181 => (x"c1",x"9a",x"c1",x"0a"),
  2182 => (x"e8",x"49",x"a2",x"c0"),
  2183 => (x"da",x"c1",x"87",x"f5"),
  2184 => (x"87",x"df",x"e6",x"49"),
  2185 => (x"d2",x"c2",x"7e",x"c1"),
  2186 => (x"66",x"c8",x"48",x"dc"),
  2187 => (x"e4",x"d2",x"c2",x"78"),
  2188 => (x"c7",x"c1",x"05",x"bf"),
  2189 => (x"c0",x"c0",x"c8",x"87"),
  2190 => (x"d0",x"d3",x"c2",x"4b"),
  2191 => (x"49",x"15",x"4d",x"7e"),
  2192 => (x"87",x"ff",x"e5",x"49"),
  2193 => (x"c0",x"02",x"98",x"70"),
  2194 => (x"b4",x"73",x"87",x"c2"),
  2195 => (x"05",x"2b",x"b7",x"c1"),
  2196 => (x"74",x"87",x"eb",x"ff"),
  2197 => (x"99",x"ff",x"c3",x"49"),
  2198 => (x"49",x"c0",x"1e",x"71"),
  2199 => (x"74",x"87",x"d1",x"fb"),
  2200 => (x"29",x"b7",x"c8",x"49"),
  2201 => (x"49",x"c1",x"1e",x"71"),
  2202 => (x"c8",x"87",x"c5",x"fb"),
  2203 => (x"49",x"fd",x"c3",x"86"),
  2204 => (x"c3",x"87",x"d0",x"e5"),
  2205 => (x"ca",x"e5",x"49",x"fa"),
  2206 => (x"87",x"fd",x"c7",x"87"),
  2207 => (x"ff",x"c3",x"49",x"74"),
  2208 => (x"2c",x"b7",x"c8",x"99"),
  2209 => (x"9c",x"74",x"b4",x"71"),
  2210 => (x"87",x"e5",x"c0",x"02"),
  2211 => (x"ff",x"48",x"a6",x"c8"),
  2212 => (x"c8",x"78",x"bf",x"c8"),
  2213 => (x"d2",x"c2",x"49",x"66"),
  2214 => (x"c2",x"89",x"bf",x"e0"),
  2215 => (x"c0",x"03",x"a9",x"e0"),
  2216 => (x"4c",x"c0",x"87",x"c5"),
  2217 => (x"c2",x"87",x"d0",x"c0"),
  2218 => (x"c8",x"48",x"e0",x"d2"),
  2219 => (x"c6",x"c0",x"78",x"66"),
  2220 => (x"e0",x"d2",x"c2",x"87"),
  2221 => (x"74",x"78",x"c0",x"48"),
  2222 => (x"05",x"99",x"c8",x"49"),
  2223 => (x"c3",x"87",x"ce",x"c0"),
  2224 => (x"fe",x"e3",x"49",x"f5"),
  2225 => (x"c2",x"49",x"70",x"87"),
  2226 => (x"e7",x"c0",x"02",x"99"),
  2227 => (x"f0",x"e6",x"c2",x"87"),
  2228 => (x"ca",x"c0",x"02",x"bf"),
  2229 => (x"88",x"c1",x"48",x"87"),
  2230 => (x"58",x"f4",x"e6",x"c2"),
  2231 => (x"c4",x"87",x"d3",x"c0"),
  2232 => (x"e0",x"c1",x"48",x"66"),
  2233 => (x"6e",x"7e",x"70",x"80"),
  2234 => (x"c5",x"c0",x"02",x"bf"),
  2235 => (x"49",x"ff",x"4b",x"87"),
  2236 => (x"7e",x"c1",x"0f",x"73"),
  2237 => (x"99",x"c4",x"49",x"74"),
  2238 => (x"87",x"ce",x"c0",x"05"),
  2239 => (x"e3",x"49",x"f2",x"c3"),
  2240 => (x"49",x"70",x"87",x"c1"),
  2241 => (x"c0",x"02",x"99",x"c2"),
  2242 => (x"e6",x"c2",x"87",x"ed"),
  2243 => (x"48",x"7e",x"bf",x"f0"),
  2244 => (x"03",x"a8",x"b7",x"c7"),
  2245 => (x"6e",x"87",x"cb",x"c0"),
  2246 => (x"c2",x"80",x"c1",x"48"),
  2247 => (x"c0",x"58",x"f4",x"e6"),
  2248 => (x"66",x"c4",x"87",x"d3"),
  2249 => (x"80",x"e0",x"c1",x"48"),
  2250 => (x"bf",x"6e",x"7e",x"70"),
  2251 => (x"87",x"c5",x"c0",x"02"),
  2252 => (x"73",x"49",x"fe",x"4b"),
  2253 => (x"c3",x"7e",x"c1",x"0f"),
  2254 => (x"c6",x"e2",x"49",x"fd"),
  2255 => (x"c2",x"49",x"70",x"87"),
  2256 => (x"e3",x"c0",x"02",x"99"),
  2257 => (x"f0",x"e6",x"c2",x"87"),
  2258 => (x"c9",x"c0",x"02",x"bf"),
  2259 => (x"f0",x"e6",x"c2",x"87"),
  2260 => (x"c0",x"78",x"c0",x"48"),
  2261 => (x"66",x"c4",x"87",x"d0"),
  2262 => (x"82",x"e0",x"c1",x"4a"),
  2263 => (x"c5",x"c0",x"02",x"6a"),
  2264 => (x"49",x"fd",x"4b",x"87"),
  2265 => (x"7e",x"c1",x"0f",x"73"),
  2266 => (x"e1",x"49",x"fa",x"c3"),
  2267 => (x"49",x"70",x"87",x"d5"),
  2268 => (x"c0",x"02",x"99",x"c2"),
  2269 => (x"e6",x"c2",x"87",x"ea"),
  2270 => (x"c7",x"48",x"bf",x"f0"),
  2271 => (x"c0",x"03",x"a8",x"b7"),
  2272 => (x"e6",x"c2",x"87",x"c9"),
  2273 => (x"78",x"c7",x"48",x"f0"),
  2274 => (x"c4",x"87",x"d3",x"c0"),
  2275 => (x"e0",x"c1",x"48",x"66"),
  2276 => (x"6e",x"7e",x"70",x"80"),
  2277 => (x"c5",x"c0",x"02",x"bf"),
  2278 => (x"49",x"fc",x"4b",x"87"),
  2279 => (x"7e",x"c1",x"0f",x"73"),
  2280 => (x"f0",x"c3",x"48",x"74"),
  2281 => (x"58",x"a6",x"cc",x"98"),
  2282 => (x"c0",x"05",x"98",x"70"),
  2283 => (x"da",x"c1",x"87",x"ce"),
  2284 => (x"87",x"cf",x"e0",x"49"),
  2285 => (x"99",x"c2",x"49",x"70"),
  2286 => (x"87",x"c1",x"c2",x"02"),
  2287 => (x"c3",x"49",x"e8",x"cf"),
  2288 => (x"a6",x"d0",x"87",x"e6"),
  2289 => (x"e8",x"e6",x"c2",x"58"),
  2290 => (x"c2",x"50",x"c0",x"48"),
  2291 => (x"bf",x"97",x"e8",x"e6"),
  2292 => (x"87",x"d9",x"c1",x"05"),
  2293 => (x"c0",x"05",x"66",x"c8"),
  2294 => (x"da",x"c1",x"87",x"cd"),
  2295 => (x"e2",x"df",x"ff",x"49"),
  2296 => (x"02",x"98",x"70",x"87"),
  2297 => (x"e8",x"87",x"c6",x"c1"),
  2298 => (x"c3",x"49",x"4b",x"bf"),
  2299 => (x"b7",x"c8",x"99",x"ff"),
  2300 => (x"c2",x"b3",x"71",x"2b"),
  2301 => (x"49",x"bf",x"e4",x"d2"),
  2302 => (x"87",x"ca",x"da",x"ff"),
  2303 => (x"c2",x"49",x"66",x"cc"),
  2304 => (x"98",x"70",x"87",x"f2"),
  2305 => (x"87",x"c6",x"c0",x"02"),
  2306 => (x"48",x"e8",x"e6",x"c2"),
  2307 => (x"e6",x"c2",x"50",x"c1"),
  2308 => (x"05",x"bf",x"97",x"e8"),
  2309 => (x"73",x"87",x"d6",x"c0"),
  2310 => (x"99",x"f0",x"c3",x"49"),
  2311 => (x"87",x"c7",x"ff",x"05"),
  2312 => (x"ff",x"49",x"da",x"c1"),
  2313 => (x"70",x"87",x"dc",x"de"),
  2314 => (x"fa",x"fe",x"05",x"98"),
  2315 => (x"f0",x"e6",x"c2",x"87"),
  2316 => (x"cc",x"4b",x"49",x"bf"),
  2317 => (x"83",x"66",x"c4",x"93"),
  2318 => (x"73",x"71",x"4b",x"6b"),
  2319 => (x"02",x"9d",x"75",x"0f"),
  2320 => (x"6d",x"87",x"e9",x"c0"),
  2321 => (x"87",x"e4",x"c0",x"02"),
  2322 => (x"dd",x"ff",x"49",x"6d"),
  2323 => (x"49",x"70",x"87",x"f5"),
  2324 => (x"c0",x"02",x"99",x"c1"),
  2325 => (x"a5",x"c4",x"87",x"cb"),
  2326 => (x"f0",x"e6",x"c2",x"4b"),
  2327 => (x"4b",x"6b",x"49",x"bf"),
  2328 => (x"02",x"85",x"c8",x"0f"),
  2329 => (x"6d",x"87",x"c5",x"c0"),
  2330 => (x"87",x"dc",x"ff",x"05"),
  2331 => (x"c8",x"c0",x"02",x"6e"),
  2332 => (x"f0",x"e6",x"c2",x"87"),
  2333 => (x"df",x"f0",x"49",x"bf"),
  2334 => (x"26",x"8e",x"f0",x"87"),
  2335 => (x"26",x"4c",x"26",x"4d"),
  2336 => (x"00",x"4f",x"26",x"4b"),
  2337 => (x"00",x"00",x"00",x"10"),
  2338 => (x"14",x"11",x"12",x"58"),
  2339 => (x"23",x"1c",x"1b",x"1d"),
  2340 => (x"94",x"91",x"59",x"5a"),
  2341 => (x"f4",x"eb",x"f2",x"f5"),
  2342 => (x"00",x"00",x"00",x"00"),
  2343 => (x"00",x"00",x"00",x"00"),
  2344 => (x"00",x"00",x"00",x"00"),
  2345 => (x"00",x"00",x"00",x"00"),
  2346 => (x"ff",x"4a",x"71",x"1e"),
  2347 => (x"72",x"49",x"bf",x"c8"),
  2348 => (x"4f",x"26",x"48",x"a1"),
  2349 => (x"bf",x"c8",x"ff",x"1e"),
  2350 => (x"c0",x"c0",x"fe",x"89"),
  2351 => (x"a9",x"c0",x"c0",x"c0"),
  2352 => (x"c0",x"87",x"c4",x"01"),
  2353 => (x"c1",x"87",x"c2",x"4a"),
  2354 => (x"26",x"48",x"72",x"4a"),
  2355 => (x"00",x"00",x"00",x"4f"),
  2356 => (x"11",x"14",x"12",x"58"),
  2357 => (x"23",x"1c",x"1b",x"1d"),
  2358 => (x"91",x"94",x"59",x"5a"),
  2359 => (x"f4",x"eb",x"f2",x"f5"),
  2360 => (x"00",x"00",x"24",x"e4"),
  2361 => (x"4f",x"54",x"55",x"41"),
  2362 => (x"54",x"4f",x"4f",x"42"),
  2363 => (x"ab",x"00",x"42",x"47"),
  2364 => (x"ab",x"00",x"00",x"19"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

